-- Custom Vendorless ROM

library ieee;
use ieee.std_logic_1164.all;

entity lane_g_root_IP is
port (
        address : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
        clock   : IN STD_LOGIC  := '1';
        q       : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
        );
end entity lane_g_root_IP;

architecture behavioral of lane_g_root_IP is
  type mem is array ( 0 to 2**12 - 1) of std_logic_vector(7 downto 0);
  constant my_Rom : mem := (
    0 => "11111111",
    1 => "11111101",
    2 => "11111011",
    3 => "11111011",
    4 => "11111010",
    5 => "11111001",
    6 => "11111001",
    7 => "11111000",
    8 => "11110111",
    9 => "11110111",
    10 => "11110111",
    11 => "11110110",
    12 => "11110110",
    13 => "11110101",
    14 => "11110101",
    15 => "11110101",
    16 => "11110100",
    17 => "11110100",
    18 => "11110011",
    19 => "11110011",
    20 => "11110011",
    21 => "11110011",
    22 => "11110010",
    23 => "11110010",
    24 => "11110010",
    25 => "11110001",
    26 => "11110001",
    27 => "11110001",
    28 => "11110001",
    29 => "11110000",
    30 => "11110000",
    31 => "11110000",
    32 => "11101111",
    33 => "11101111",
    34 => "11101111",
    35 => "11101111",
    36 => "11101111",
    37 => "11101110",
    38 => "11101110",
    39 => "11101110",
    40 => "11101110",
    41 => "11101101",
    42 => "11101101",
    43 => "11101101",
    44 => "11101101",
    45 => "11101101",
    46 => "11101100",
    47 => "11101100",
    48 => "11101100",
    49 => "11101100",
    50 => "11101011",
    51 => "11101011",
    52 => "11101011",
    53 => "11101011",
    54 => "11101011",
    55 => "11101011",
    56 => "11101010",
    57 => "11101010",
    58 => "11101010",
    59 => "11101010",
    60 => "11101010",
    61 => "11101001",
    62 => "11101001",
    63 => "11101001",
    64 => "11101001",
    65 => "11101001",
    66 => "11101001",
    67 => "11101000",
    68 => "11101000",
    69 => "11101000",
    70 => "11101000",
    71 => "11101000",
    72 => "11100111",
    73 => "11100111",
    74 => "11100111",
    75 => "11100111",
    76 => "11100111",
    77 => "11100111",
    78 => "11100111",
    79 => "11100110",
    80 => "11100110",
    81 => "11100110",
    82 => "11100110",
    83 => "11100110",
    84 => "11100110",
    85 => "11100101",
    86 => "11100101",
    87 => "11100101",
    88 => "11100101",
    89 => "11100101",
    90 => "11100101",
    91 => "11100101",
    92 => "11100100",
    93 => "11100100",
    94 => "11100100",
    95 => "11100100",
    96 => "11100100",
    97 => "11100100",
    98 => "11100011",
    99 => "11100011",
    100 => "11100011",
    101 => "11100011",
    102 => "11100011",
    103 => "11100011",
    104 => "11100011",
    105 => "11100011",
    106 => "11100010",
    107 => "11100010",
    108 => "11100010",
    109 => "11100010",
    110 => "11100010",
    111 => "11100010",
    112 => "11100010",
    113 => "11100001",
    114 => "11100001",
    115 => "11100001",
    116 => "11100001",
    117 => "11100001",
    118 => "11100001",
    119 => "11100001",
    120 => "11100001",
    121 => "11100000",
    122 => "11100000",
    123 => "11100000",
    124 => "11100000",
    125 => "11100000",
    126 => "11100000",
    127 => "11100000",
    128 => "11011111",
    129 => "11011111",
    130 => "11011111",
    131 => "11011111",
    132 => "11011111",
    133 => "11011111",
    134 => "11011111",
    135 => "11011111",
    136 => "11011111",
    137 => "11011110",
    138 => "11011110",
    139 => "11011110",
    140 => "11011110",
    141 => "11011110",
    142 => "11011110",
    143 => "11011110",
    144 => "11011110",
    145 => "11011101",
    146 => "11011101",
    147 => "11011101",
    148 => "11011101",
    149 => "11011101",
    150 => "11011101",
    151 => "11011101",
    152 => "11011101",
    153 => "11011101",
    154 => "11011100",
    155 => "11011100",
    156 => "11011100",
    157 => "11011100",
    158 => "11011100",
    159 => "11011100",
    160 => "11011100",
    161 => "11011100",
    162 => "11011011",
    163 => "11011011",
    164 => "11011011",
    165 => "11011011",
    166 => "11011011",
    167 => "11011011",
    168 => "11011011",
    169 => "11011011",
    170 => "11011011",
    171 => "11011011",
    172 => "11011010",
    173 => "11011010",
    174 => "11011010",
    175 => "11011010",
    176 => "11011010",
    177 => "11011010",
    178 => "11011010",
    179 => "11011010",
    180 => "11011010",
    181 => "11011001",
    182 => "11011001",
    183 => "11011001",
    184 => "11011001",
    185 => "11011001",
    186 => "11011001",
    187 => "11011001",
    188 => "11011001",
    189 => "11011001",
    190 => "11011001",
    191 => "11011000",
    192 => "11011000",
    193 => "11011000",
    194 => "11011000",
    195 => "11011000",
    196 => "11011000",
    197 => "11011000",
    198 => "11011000",
    199 => "11011000",
    200 => "11010111",
    201 => "11010111",
    202 => "11010111",
    203 => "11010111",
    204 => "11010111",
    205 => "11010111",
    206 => "11010111",
    207 => "11010111",
    208 => "11010111",
    209 => "11010111",
    210 => "11010111",
    211 => "11010110",
    212 => "11010110",
    213 => "11010110",
    214 => "11010110",
    215 => "11010110",
    216 => "11010110",
    217 => "11010110",
    218 => "11010110",
    219 => "11010110",
    220 => "11010110",
    221 => "11010101",
    222 => "11010101",
    223 => "11010101",
    224 => "11010101",
    225 => "11010101",
    226 => "11010101",
    227 => "11010101",
    228 => "11010101",
    229 => "11010101",
    230 => "11010101",
    231 => "11010101",
    232 => "11010100",
    233 => "11010100",
    234 => "11010100",
    235 => "11010100",
    236 => "11010100",
    237 => "11010100",
    238 => "11010100",
    239 => "11010100",
    240 => "11010100",
    241 => "11010100",
    242 => "11010011",
    243 => "11010011",
    244 => "11010011",
    245 => "11010011",
    246 => "11010011",
    247 => "11010011",
    248 => "11010011",
    249 => "11010011",
    250 => "11010011",
    251 => "11010011",
    252 => "11010011",
    253 => "11010011",
    254 => "11010010",
    255 => "11010010",
    256 => "11010010",
    257 => "11010010",
    258 => "11010010",
    259 => "11010010",
    260 => "11010010",
    261 => "11010010",
    262 => "11010010",
    263 => "11010010",
    264 => "11010010",
    265 => "11010001",
    266 => "11010001",
    267 => "11010001",
    268 => "11010001",
    269 => "11010001",
    270 => "11010001",
    271 => "11010001",
    272 => "11010001",
    273 => "11010001",
    274 => "11010001",
    275 => "11010001",
    276 => "11010001",
    277 => "11010000",
    278 => "11010000",
    279 => "11010000",
    280 => "11010000",
    281 => "11010000",
    282 => "11010000",
    283 => "11010000",
    284 => "11010000",
    285 => "11010000",
    286 => "11010000",
    287 => "11010000",
    288 => "11001111",
    289 => "11001111",
    290 => "11001111",
    291 => "11001111",
    292 => "11001111",
    293 => "11001111",
    294 => "11001111",
    295 => "11001111",
    296 => "11001111",
    297 => "11001111",
    298 => "11001111",
    299 => "11001111",
    300 => "11001111",
    301 => "11001110",
    302 => "11001110",
    303 => "11001110",
    304 => "11001110",
    305 => "11001110",
    306 => "11001110",
    307 => "11001110",
    308 => "11001110",
    309 => "11001110",
    310 => "11001110",
    311 => "11001110",
    312 => "11001110",
    313 => "11001101",
    314 => "11001101",
    315 => "11001101",
    316 => "11001101",
    317 => "11001101",
    318 => "11001101",
    319 => "11001101",
    320 => "11001101",
    321 => "11001101",
    322 => "11001101",
    323 => "11001101",
    324 => "11001101",
    325 => "11001101",
    326 => "11001100",
    327 => "11001100",
    328 => "11001100",
    329 => "11001100",
    330 => "11001100",
    331 => "11001100",
    332 => "11001100",
    333 => "11001100",
    334 => "11001100",
    335 => "11001100",
    336 => "11001100",
    337 => "11001100",
    338 => "11001011",
    339 => "11001011",
    340 => "11001011",
    341 => "11001011",
    342 => "11001011",
    343 => "11001011",
    344 => "11001011",
    345 => "11001011",
    346 => "11001011",
    347 => "11001011",
    348 => "11001011",
    349 => "11001011",
    350 => "11001011",
    351 => "11001011",
    352 => "11001010",
    353 => "11001010",
    354 => "11001010",
    355 => "11001010",
    356 => "11001010",
    357 => "11001010",
    358 => "11001010",
    359 => "11001010",
    360 => "11001010",
    361 => "11001010",
    362 => "11001010",
    363 => "11001010",
    364 => "11001010",
    365 => "11001001",
    366 => "11001001",
    367 => "11001001",
    368 => "11001001",
    369 => "11001001",
    370 => "11001001",
    371 => "11001001",
    372 => "11001001",
    373 => "11001001",
    374 => "11001001",
    375 => "11001001",
    376 => "11001001",
    377 => "11001001",
    378 => "11001001",
    379 => "11001000",
    380 => "11001000",
    381 => "11001000",
    382 => "11001000",
    383 => "11001000",
    384 => "11001000",
    385 => "11001000",
    386 => "11001000",
    387 => "11001000",
    388 => "11001000",
    389 => "11001000",
    390 => "11001000",
    391 => "11001000",
    392 => "11000111",
    393 => "11000111",
    394 => "11000111",
    395 => "11000111",
    396 => "11000111",
    397 => "11000111",
    398 => "11000111",
    399 => "11000111",
    400 => "11000111",
    401 => "11000111",
    402 => "11000111",
    403 => "11000111",
    404 => "11000111",
    405 => "11000111",
    406 => "11000111",
    407 => "11000110",
    408 => "11000110",
    409 => "11000110",
    410 => "11000110",
    411 => "11000110",
    412 => "11000110",
    413 => "11000110",
    414 => "11000110",
    415 => "11000110",
    416 => "11000110",
    417 => "11000110",
    418 => "11000110",
    419 => "11000110",
    420 => "11000110",
    421 => "11000101",
    422 => "11000101",
    423 => "11000101",
    424 => "11000101",
    425 => "11000101",
    426 => "11000101",
    427 => "11000101",
    428 => "11000101",
    429 => "11000101",
    430 => "11000101",
    431 => "11000101",
    432 => "11000101",
    433 => "11000101",
    434 => "11000101",
    435 => "11000101",
    436 => "11000100",
    437 => "11000100",
    438 => "11000100",
    439 => "11000100",
    440 => "11000100",
    441 => "11000100",
    442 => "11000100",
    443 => "11000100",
    444 => "11000100",
    445 => "11000100",
    446 => "11000100",
    447 => "11000100",
    448 => "11000100",
    449 => "11000100",
    450 => "11000011",
    451 => "11000011",
    452 => "11000011",
    453 => "11000011",
    454 => "11000011",
    455 => "11000011",
    456 => "11000011",
    457 => "11000011",
    458 => "11000011",
    459 => "11000011",
    460 => "11000011",
    461 => "11000011",
    462 => "11000011",
    463 => "11000011",
    464 => "11000011",
    465 => "11000011",
    466 => "11000010",
    467 => "11000010",
    468 => "11000010",
    469 => "11000010",
    470 => "11000010",
    471 => "11000010",
    472 => "11000010",
    473 => "11000010",
    474 => "11000010",
    475 => "11000010",
    476 => "11000010",
    477 => "11000010",
    478 => "11000010",
    479 => "11000010",
    480 => "11000010",
    481 => "11000001",
    482 => "11000001",
    483 => "11000001",
    484 => "11000001",
    485 => "11000001",
    486 => "11000001",
    487 => "11000001",
    488 => "11000001",
    489 => "11000001",
    490 => "11000001",
    491 => "11000001",
    492 => "11000001",
    493 => "11000001",
    494 => "11000001",
    495 => "11000001",
    496 => "11000001",
    497 => "11000000",
    498 => "11000000",
    499 => "11000000",
    500 => "11000000",
    501 => "11000000",
    502 => "11000000",
    503 => "11000000",
    504 => "11000000",
    505 => "11000000",
    506 => "11000000",
    507 => "11000000",
    508 => "11000000",
    509 => "11000000",
    510 => "11000000",
    511 => "11000000",
    512 => "10111111",
    513 => "10111111",
    514 => "10111111",
    515 => "10111111",
    516 => "10111111",
    517 => "10111111",
    518 => "10111111",
    519 => "10111111",
    520 => "10111111",
    521 => "10111111",
    522 => "10111111",
    523 => "10111111",
    524 => "10111111",
    525 => "10111111",
    526 => "10111111",
    527 => "10111111",
    528 => "10111111",
    529 => "10111110",
    530 => "10111110",
    531 => "10111110",
    532 => "10111110",
    533 => "10111110",
    534 => "10111110",
    535 => "10111110",
    536 => "10111110",
    537 => "10111110",
    538 => "10111110",
    539 => "10111110",
    540 => "10111110",
    541 => "10111110",
    542 => "10111110",
    543 => "10111110",
    544 => "10111110",
    545 => "10111101",
    546 => "10111101",
    547 => "10111101",
    548 => "10111101",
    549 => "10111101",
    550 => "10111101",
    551 => "10111101",
    552 => "10111101",
    553 => "10111101",
    554 => "10111101",
    555 => "10111101",
    556 => "10111101",
    557 => "10111101",
    558 => "10111101",
    559 => "10111101",
    560 => "10111101",
    561 => "10111101",
    562 => "10111100",
    563 => "10111100",
    564 => "10111100",
    565 => "10111100",
    566 => "10111100",
    567 => "10111100",
    568 => "10111100",
    569 => "10111100",
    570 => "10111100",
    571 => "10111100",
    572 => "10111100",
    573 => "10111100",
    574 => "10111100",
    575 => "10111100",
    576 => "10111100",
    577 => "10111100",
    578 => "10111011",
    579 => "10111011",
    580 => "10111011",
    581 => "10111011",
    582 => "10111011",
    583 => "10111011",
    584 => "10111011",
    585 => "10111011",
    586 => "10111011",
    587 => "10111011",
    588 => "10111011",
    589 => "10111011",
    590 => "10111011",
    591 => "10111011",
    592 => "10111011",
    593 => "10111011",
    594 => "10111011",
    595 => "10111011",
    596 => "10111010",
    597 => "10111010",
    598 => "10111010",
    599 => "10111010",
    600 => "10111010",
    601 => "10111010",
    602 => "10111010",
    603 => "10111010",
    604 => "10111010",
    605 => "10111010",
    606 => "10111010",
    607 => "10111010",
    608 => "10111010",
    609 => "10111010",
    610 => "10111010",
    611 => "10111010",
    612 => "10111010",
    613 => "10111001",
    614 => "10111001",
    615 => "10111001",
    616 => "10111001",
    617 => "10111001",
    618 => "10111001",
    619 => "10111001",
    620 => "10111001",
    621 => "10111001",
    622 => "10111001",
    623 => "10111001",
    624 => "10111001",
    625 => "10111001",
    626 => "10111001",
    627 => "10111001",
    628 => "10111001",
    629 => "10111001",
    630 => "10111001",
    631 => "10111000",
    632 => "10111000",
    633 => "10111000",
    634 => "10111000",
    635 => "10111000",
    636 => "10111000",
    637 => "10111000",
    638 => "10111000",
    639 => "10111000",
    640 => "10111000",
    641 => "10111000",
    642 => "10111000",
    643 => "10111000",
    644 => "10111000",
    645 => "10111000",
    646 => "10111000",
    647 => "10111000",
    648 => "10110111",
    649 => "10110111",
    650 => "10110111",
    651 => "10110111",
    652 => "10110111",
    653 => "10110111",
    654 => "10110111",
    655 => "10110111",
    656 => "10110111",
    657 => "10110111",
    658 => "10110111",
    659 => "10110111",
    660 => "10110111",
    661 => "10110111",
    662 => "10110111",
    663 => "10110111",
    664 => "10110111",
    665 => "10110111",
    666 => "10110111",
    667 => "10110110",
    668 => "10110110",
    669 => "10110110",
    670 => "10110110",
    671 => "10110110",
    672 => "10110110",
    673 => "10110110",
    674 => "10110110",
    675 => "10110110",
    676 => "10110110",
    677 => "10110110",
    678 => "10110110",
    679 => "10110110",
    680 => "10110110",
    681 => "10110110",
    682 => "10110110",
    683 => "10110110",
    684 => "10110110",
    685 => "10110101",
    686 => "10110101",
    687 => "10110101",
    688 => "10110101",
    689 => "10110101",
    690 => "10110101",
    691 => "10110101",
    692 => "10110101",
    693 => "10110101",
    694 => "10110101",
    695 => "10110101",
    696 => "10110101",
    697 => "10110101",
    698 => "10110101",
    699 => "10110101",
    700 => "10110101",
    701 => "10110101",
    702 => "10110101",
    703 => "10110101",
    704 => "10110100",
    705 => "10110100",
    706 => "10110100",
    707 => "10110100",
    708 => "10110100",
    709 => "10110100",
    710 => "10110100",
    711 => "10110100",
    712 => "10110100",
    713 => "10110100",
    714 => "10110100",
    715 => "10110100",
    716 => "10110100",
    717 => "10110100",
    718 => "10110100",
    719 => "10110100",
    720 => "10110100",
    721 => "10110100",
    722 => "10110011",
    723 => "10110011",
    724 => "10110011",
    725 => "10110011",
    726 => "10110011",
    727 => "10110011",
    728 => "10110011",
    729 => "10110011",
    730 => "10110011",
    731 => "10110011",
    732 => "10110011",
    733 => "10110011",
    734 => "10110011",
    735 => "10110011",
    736 => "10110011",
    737 => "10110011",
    738 => "10110011",
    739 => "10110011",
    740 => "10110011",
    741 => "10110011",
    742 => "10110010",
    743 => "10110010",
    744 => "10110010",
    745 => "10110010",
    746 => "10110010",
    747 => "10110010",
    748 => "10110010",
    749 => "10110010",
    750 => "10110010",
    751 => "10110010",
    752 => "10110010",
    753 => "10110010",
    754 => "10110010",
    755 => "10110010",
    756 => "10110010",
    757 => "10110010",
    758 => "10110010",
    759 => "10110010",
    760 => "10110010",
    761 => "10110001",
    762 => "10110001",
    763 => "10110001",
    764 => "10110001",
    765 => "10110001",
    766 => "10110001",
    767 => "10110001",
    768 => "10110001",
    769 => "10110001",
    770 => "10110001",
    771 => "10110001",
    772 => "10110001",
    773 => "10110001",
    774 => "10110001",
    775 => "10110001",
    776 => "10110001",
    777 => "10110001",
    778 => "10110001",
    779 => "10110001",
    780 => "10110001",
    781 => "10110000",
    782 => "10110000",
    783 => "10110000",
    784 => "10110000",
    785 => "10110000",
    786 => "10110000",
    787 => "10110000",
    788 => "10110000",
    789 => "10110000",
    790 => "10110000",
    791 => "10110000",
    792 => "10110000",
    793 => "10110000",
    794 => "10110000",
    795 => "10110000",
    796 => "10110000",
    797 => "10110000",
    798 => "10110000",
    799 => "10110000",
    800 => "10101111",
    801 => "10101111",
    802 => "10101111",
    803 => "10101111",
    804 => "10101111",
    805 => "10101111",
    806 => "10101111",
    807 => "10101111",
    808 => "10101111",
    809 => "10101111",
    810 => "10101111",
    811 => "10101111",
    812 => "10101111",
    813 => "10101111",
    814 => "10101111",
    815 => "10101111",
    816 => "10101111",
    817 => "10101111",
    818 => "10101111",
    819 => "10101111",
    820 => "10101111",
    821 => "10101110",
    822 => "10101110",
    823 => "10101110",
    824 => "10101110",
    825 => "10101110",
    826 => "10101110",
    827 => "10101110",
    828 => "10101110",
    829 => "10101110",
    830 => "10101110",
    831 => "10101110",
    832 => "10101110",
    833 => "10101110",
    834 => "10101110",
    835 => "10101110",
    836 => "10101110",
    837 => "10101110",
    838 => "10101110",
    839 => "10101110",
    840 => "10101110",
    841 => "10101101",
    842 => "10101101",
    843 => "10101101",
    844 => "10101101",
    845 => "10101101",
    846 => "10101101",
    847 => "10101101",
    848 => "10101101",
    849 => "10101101",
    850 => "10101101",
    851 => "10101101",
    852 => "10101101",
    853 => "10101101",
    854 => "10101101",
    855 => "10101101",
    856 => "10101101",
    857 => "10101101",
    858 => "10101101",
    859 => "10101101",
    860 => "10101101",
    861 => "10101101",
    862 => "10101100",
    863 => "10101100",
    864 => "10101100",
    865 => "10101100",
    866 => "10101100",
    867 => "10101100",
    868 => "10101100",
    869 => "10101100",
    870 => "10101100",
    871 => "10101100",
    872 => "10101100",
    873 => "10101100",
    874 => "10101100",
    875 => "10101100",
    876 => "10101100",
    877 => "10101100",
    878 => "10101100",
    879 => "10101100",
    880 => "10101100",
    881 => "10101100",
    882 => "10101011",
    883 => "10101011",
    884 => "10101011",
    885 => "10101011",
    886 => "10101011",
    887 => "10101011",
    888 => "10101011",
    889 => "10101011",
    890 => "10101011",
    891 => "10101011",
    892 => "10101011",
    893 => "10101011",
    894 => "10101011",
    895 => "10101011",
    896 => "10101011",
    897 => "10101011",
    898 => "10101011",
    899 => "10101011",
    900 => "10101011",
    901 => "10101011",
    902 => "10101011",
    903 => "10101011",
    904 => "10101010",
    905 => "10101010",
    906 => "10101010",
    907 => "10101010",
    908 => "10101010",
    909 => "10101010",
    910 => "10101010",
    911 => "10101010",
    912 => "10101010",
    913 => "10101010",
    914 => "10101010",
    915 => "10101010",
    916 => "10101010",
    917 => "10101010",
    918 => "10101010",
    919 => "10101010",
    920 => "10101010",
    921 => "10101010",
    922 => "10101010",
    923 => "10101010",
    924 => "10101010",
    925 => "10101001",
    926 => "10101001",
    927 => "10101001",
    928 => "10101001",
    929 => "10101001",
    930 => "10101001",
    931 => "10101001",
    932 => "10101001",
    933 => "10101001",
    934 => "10101001",
    935 => "10101001",
    936 => "10101001",
    937 => "10101001",
    938 => "10101001",
    939 => "10101001",
    940 => "10101001",
    941 => "10101001",
    942 => "10101001",
    943 => "10101001",
    944 => "10101001",
    945 => "10101001",
    946 => "10101001",
    947 => "10101000",
    948 => "10101000",
    949 => "10101000",
    950 => "10101000",
    951 => "10101000",
    952 => "10101000",
    953 => "10101000",
    954 => "10101000",
    955 => "10101000",
    956 => "10101000",
    957 => "10101000",
    958 => "10101000",
    959 => "10101000",
    960 => "10101000",
    961 => "10101000",
    962 => "10101000",
    963 => "10101000",
    964 => "10101000",
    965 => "10101000",
    966 => "10101000",
    967 => "10101000",
    968 => "10100111",
    969 => "10100111",
    970 => "10100111",
    971 => "10100111",
    972 => "10100111",
    973 => "10100111",
    974 => "10100111",
    975 => "10100111",
    976 => "10100111",
    977 => "10100111",
    978 => "10100111",
    979 => "10100111",
    980 => "10100111",
    981 => "10100111",
    982 => "10100111",
    983 => "10100111",
    984 => "10100111",
    985 => "10100111",
    986 => "10100111",
    987 => "10100111",
    988 => "10100111",
    989 => "10100111",
    990 => "10100111",
    991 => "10100110",
    992 => "10100110",
    993 => "10100110",
    994 => "10100110",
    995 => "10100110",
    996 => "10100110",
    997 => "10100110",
    998 => "10100110",
    999 => "10100110",
    1000 => "10100110",
    1001 => "10100110",
    1002 => "10100110",
    1003 => "10100110",
    1004 => "10100110",
    1005 => "10100110",
    1006 => "10100110",
    1007 => "10100110",
    1008 => "10100110",
    1009 => "10100110",
    1010 => "10100110",
    1011 => "10100110",
    1012 => "10100110",
    1013 => "10100101",
    1014 => "10100101",
    1015 => "10100101",
    1016 => "10100101",
    1017 => "10100101",
    1018 => "10100101",
    1019 => "10100101",
    1020 => "10100101",
    1021 => "10100101",
    1022 => "10100101",
    1023 => "10100101",
    1024 => "10100101",
    1025 => "10100101",
    1026 => "10100101",
    1027 => "10100101",
    1028 => "10100101",
    1029 => "10100101",
    1030 => "10100101",
    1031 => "10100101",
    1032 => "10100101",
    1033 => "10100101",
    1034 => "10100101",
    1035 => "10100101",
    1036 => "10100100",
    1037 => "10100100",
    1038 => "10100100",
    1039 => "10100100",
    1040 => "10100100",
    1041 => "10100100",
    1042 => "10100100",
    1043 => "10100100",
    1044 => "10100100",
    1045 => "10100100",
    1046 => "10100100",
    1047 => "10100100",
    1048 => "10100100",
    1049 => "10100100",
    1050 => "10100100",
    1051 => "10100100",
    1052 => "10100100",
    1053 => "10100100",
    1054 => "10100100",
    1055 => "10100100",
    1056 => "10100100",
    1057 => "10100100",
    1058 => "10100011",
    1059 => "10100011",
    1060 => "10100011",
    1061 => "10100011",
    1062 => "10100011",
    1063 => "10100011",
    1064 => "10100011",
    1065 => "10100011",
    1066 => "10100011",
    1067 => "10100011",
    1068 => "10100011",
    1069 => "10100011",
    1070 => "10100011",
    1071 => "10100011",
    1072 => "10100011",
    1073 => "10100011",
    1074 => "10100011",
    1075 => "10100011",
    1076 => "10100011",
    1077 => "10100011",
    1078 => "10100011",
    1079 => "10100011",
    1080 => "10100011",
    1081 => "10100011",
    1082 => "10100010",
    1083 => "10100010",
    1084 => "10100010",
    1085 => "10100010",
    1086 => "10100010",
    1087 => "10100010",
    1088 => "10100010",
    1089 => "10100010",
    1090 => "10100010",
    1091 => "10100010",
    1092 => "10100010",
    1093 => "10100010",
    1094 => "10100010",
    1095 => "10100010",
    1096 => "10100010",
    1097 => "10100010",
    1098 => "10100010",
    1099 => "10100010",
    1100 => "10100010",
    1101 => "10100010",
    1102 => "10100010",
    1103 => "10100010",
    1104 => "10100010",
    1105 => "10100001",
    1106 => "10100001",
    1107 => "10100001",
    1108 => "10100001",
    1109 => "10100001",
    1110 => "10100001",
    1111 => "10100001",
    1112 => "10100001",
    1113 => "10100001",
    1114 => "10100001",
    1115 => "10100001",
    1116 => "10100001",
    1117 => "10100001",
    1118 => "10100001",
    1119 => "10100001",
    1120 => "10100001",
    1121 => "10100001",
    1122 => "10100001",
    1123 => "10100001",
    1124 => "10100001",
    1125 => "10100001",
    1126 => "10100001",
    1127 => "10100001",
    1128 => "10100001",
    1129 => "10100000",
    1130 => "10100000",
    1131 => "10100000",
    1132 => "10100000",
    1133 => "10100000",
    1134 => "10100000",
    1135 => "10100000",
    1136 => "10100000",
    1137 => "10100000",
    1138 => "10100000",
    1139 => "10100000",
    1140 => "10100000",
    1141 => "10100000",
    1142 => "10100000",
    1143 => "10100000",
    1144 => "10100000",
    1145 => "10100000",
    1146 => "10100000",
    1147 => "10100000",
    1148 => "10100000",
    1149 => "10100000",
    1150 => "10100000",
    1151 => "10100000",
    1152 => "10011111",
    1153 => "10011111",
    1154 => "10011111",
    1155 => "10011111",
    1156 => "10011111",
    1157 => "10011111",
    1158 => "10011111",
    1159 => "10011111",
    1160 => "10011111",
    1161 => "10011111",
    1162 => "10011111",
    1163 => "10011111",
    1164 => "10011111",
    1165 => "10011111",
    1166 => "10011111",
    1167 => "10011111",
    1168 => "10011111",
    1169 => "10011111",
    1170 => "10011111",
    1171 => "10011111",
    1172 => "10011111",
    1173 => "10011111",
    1174 => "10011111",
    1175 => "10011111",
    1176 => "10011111",
    1177 => "10011110",
    1178 => "10011110",
    1179 => "10011110",
    1180 => "10011110",
    1181 => "10011110",
    1182 => "10011110",
    1183 => "10011110",
    1184 => "10011110",
    1185 => "10011110",
    1186 => "10011110",
    1187 => "10011110",
    1188 => "10011110",
    1189 => "10011110",
    1190 => "10011110",
    1191 => "10011110",
    1192 => "10011110",
    1193 => "10011110",
    1194 => "10011110",
    1195 => "10011110",
    1196 => "10011110",
    1197 => "10011110",
    1198 => "10011110",
    1199 => "10011110",
    1200 => "10011110",
    1201 => "10011101",
    1202 => "10011101",
    1203 => "10011101",
    1204 => "10011101",
    1205 => "10011101",
    1206 => "10011101",
    1207 => "10011101",
    1208 => "10011101",
    1209 => "10011101",
    1210 => "10011101",
    1211 => "10011101",
    1212 => "10011101",
    1213 => "10011101",
    1214 => "10011101",
    1215 => "10011101",
    1216 => "10011101",
    1217 => "10011101",
    1218 => "10011101",
    1219 => "10011101",
    1220 => "10011101",
    1221 => "10011101",
    1222 => "10011101",
    1223 => "10011101",
    1224 => "10011101",
    1225 => "10011101",
    1226 => "10011100",
    1227 => "10011100",
    1228 => "10011100",
    1229 => "10011100",
    1230 => "10011100",
    1231 => "10011100",
    1232 => "10011100",
    1233 => "10011100",
    1234 => "10011100",
    1235 => "10011100",
    1236 => "10011100",
    1237 => "10011100",
    1238 => "10011100",
    1239 => "10011100",
    1240 => "10011100",
    1241 => "10011100",
    1242 => "10011100",
    1243 => "10011100",
    1244 => "10011100",
    1245 => "10011100",
    1246 => "10011100",
    1247 => "10011100",
    1248 => "10011100",
    1249 => "10011100",
    1250 => "10011011",
    1251 => "10011011",
    1252 => "10011011",
    1253 => "10011011",
    1254 => "10011011",
    1255 => "10011011",
    1256 => "10011011",
    1257 => "10011011",
    1258 => "10011011",
    1259 => "10011011",
    1260 => "10011011",
    1261 => "10011011",
    1262 => "10011011",
    1263 => "10011011",
    1264 => "10011011",
    1265 => "10011011",
    1266 => "10011011",
    1267 => "10011011",
    1268 => "10011011",
    1269 => "10011011",
    1270 => "10011011",
    1271 => "10011011",
    1272 => "10011011",
    1273 => "10011011",
    1274 => "10011011",
    1275 => "10011011",
    1276 => "10011010",
    1277 => "10011010",
    1278 => "10011010",
    1279 => "10011010",
    1280 => "10011010",
    1281 => "10011010",
    1282 => "10011010",
    1283 => "10011010",
    1284 => "10011010",
    1285 => "10011010",
    1286 => "10011010",
    1287 => "10011010",
    1288 => "10011010",
    1289 => "10011010",
    1290 => "10011010",
    1291 => "10011010",
    1292 => "10011010",
    1293 => "10011010",
    1294 => "10011010",
    1295 => "10011010",
    1296 => "10011010",
    1297 => "10011010",
    1298 => "10011010",
    1299 => "10011010",
    1300 => "10011010",
    1301 => "10011001",
    1302 => "10011001",
    1303 => "10011001",
    1304 => "10011001",
    1305 => "10011001",
    1306 => "10011001",
    1307 => "10011001",
    1308 => "10011001",
    1309 => "10011001",
    1310 => "10011001",
    1311 => "10011001",
    1312 => "10011001",
    1313 => "10011001",
    1314 => "10011001",
    1315 => "10011001",
    1316 => "10011001",
    1317 => "10011001",
    1318 => "10011001",
    1319 => "10011001",
    1320 => "10011001",
    1321 => "10011001",
    1322 => "10011001",
    1323 => "10011001",
    1324 => "10011001",
    1325 => "10011001",
    1326 => "10011001",
    1327 => "10011000",
    1328 => "10011000",
    1329 => "10011000",
    1330 => "10011000",
    1331 => "10011000",
    1332 => "10011000",
    1333 => "10011000",
    1334 => "10011000",
    1335 => "10011000",
    1336 => "10011000",
    1337 => "10011000",
    1338 => "10011000",
    1339 => "10011000",
    1340 => "10011000",
    1341 => "10011000",
    1342 => "10011000",
    1343 => "10011000",
    1344 => "10011000",
    1345 => "10011000",
    1346 => "10011000",
    1347 => "10011000",
    1348 => "10011000",
    1349 => "10011000",
    1350 => "10011000",
    1351 => "10011000",
    1352 => "10010111",
    1353 => "10010111",
    1354 => "10010111",
    1355 => "10010111",
    1356 => "10010111",
    1357 => "10010111",
    1358 => "10010111",
    1359 => "10010111",
    1360 => "10010111",
    1361 => "10010111",
    1362 => "10010111",
    1363 => "10010111",
    1364 => "10010111",
    1365 => "10010111",
    1366 => "10010111",
    1367 => "10010111",
    1368 => "10010111",
    1369 => "10010111",
    1370 => "10010111",
    1371 => "10010111",
    1372 => "10010111",
    1373 => "10010111",
    1374 => "10010111",
    1375 => "10010111",
    1376 => "10010111",
    1377 => "10010111",
    1378 => "10010111",
    1379 => "10010110",
    1380 => "10010110",
    1381 => "10010110",
    1382 => "10010110",
    1383 => "10010110",
    1384 => "10010110",
    1385 => "10010110",
    1386 => "10010110",
    1387 => "10010110",
    1388 => "10010110",
    1389 => "10010110",
    1390 => "10010110",
    1391 => "10010110",
    1392 => "10010110",
    1393 => "10010110",
    1394 => "10010110",
    1395 => "10010110",
    1396 => "10010110",
    1397 => "10010110",
    1398 => "10010110",
    1399 => "10010110",
    1400 => "10010110",
    1401 => "10010110",
    1402 => "10010110",
    1403 => "10010110",
    1404 => "10010110",
    1405 => "10010101",
    1406 => "10010101",
    1407 => "10010101",
    1408 => "10010101",
    1409 => "10010101",
    1410 => "10010101",
    1411 => "10010101",
    1412 => "10010101",
    1413 => "10010101",
    1414 => "10010101",
    1415 => "10010101",
    1416 => "10010101",
    1417 => "10010101",
    1418 => "10010101",
    1419 => "10010101",
    1420 => "10010101",
    1421 => "10010101",
    1422 => "10010101",
    1423 => "10010101",
    1424 => "10010101",
    1425 => "10010101",
    1426 => "10010101",
    1427 => "10010101",
    1428 => "10010101",
    1429 => "10010101",
    1430 => "10010101",
    1431 => "10010101",
    1432 => "10010100",
    1433 => "10010100",
    1434 => "10010100",
    1435 => "10010100",
    1436 => "10010100",
    1437 => "10010100",
    1438 => "10010100",
    1439 => "10010100",
    1440 => "10010100",
    1441 => "10010100",
    1442 => "10010100",
    1443 => "10010100",
    1444 => "10010100",
    1445 => "10010100",
    1446 => "10010100",
    1447 => "10010100",
    1448 => "10010100",
    1449 => "10010100",
    1450 => "10010100",
    1451 => "10010100",
    1452 => "10010100",
    1453 => "10010100",
    1454 => "10010100",
    1455 => "10010100",
    1456 => "10010100",
    1457 => "10010100",
    1458 => "10010011",
    1459 => "10010011",
    1460 => "10010011",
    1461 => "10010011",
    1462 => "10010011",
    1463 => "10010011",
    1464 => "10010011",
    1465 => "10010011",
    1466 => "10010011",
    1467 => "10010011",
    1468 => "10010011",
    1469 => "10010011",
    1470 => "10010011",
    1471 => "10010011",
    1472 => "10010011",
    1473 => "10010011",
    1474 => "10010011",
    1475 => "10010011",
    1476 => "10010011",
    1477 => "10010011",
    1478 => "10010011",
    1479 => "10010011",
    1480 => "10010011",
    1481 => "10010011",
    1482 => "10010011",
    1483 => "10010011",
    1484 => "10010011",
    1485 => "10010011",
    1486 => "10010010",
    1487 => "10010010",
    1488 => "10010010",
    1489 => "10010010",
    1490 => "10010010",
    1491 => "10010010",
    1492 => "10010010",
    1493 => "10010010",
    1494 => "10010010",
    1495 => "10010010",
    1496 => "10010010",
    1497 => "10010010",
    1498 => "10010010",
    1499 => "10010010",
    1500 => "10010010",
    1501 => "10010010",
    1502 => "10010010",
    1503 => "10010010",
    1504 => "10010010",
    1505 => "10010010",
    1506 => "10010010",
    1507 => "10010010",
    1508 => "10010010",
    1509 => "10010010",
    1510 => "10010010",
    1511 => "10010010",
    1512 => "10010010",
    1513 => "10010001",
    1514 => "10010001",
    1515 => "10010001",
    1516 => "10010001",
    1517 => "10010001",
    1518 => "10010001",
    1519 => "10010001",
    1520 => "10010001",
    1521 => "10010001",
    1522 => "10010001",
    1523 => "10010001",
    1524 => "10010001",
    1525 => "10010001",
    1526 => "10010001",
    1527 => "10010001",
    1528 => "10010001",
    1529 => "10010001",
    1530 => "10010001",
    1531 => "10010001",
    1532 => "10010001",
    1533 => "10010001",
    1534 => "10010001",
    1535 => "10010001",
    1536 => "10010001",
    1537 => "10010001",
    1538 => "10010001",
    1539 => "10010001",
    1540 => "10010001",
    1541 => "10010000",
    1542 => "10010000",
    1543 => "10010000",
    1544 => "10010000",
    1545 => "10010000",
    1546 => "10010000",
    1547 => "10010000",
    1548 => "10010000",
    1549 => "10010000",
    1550 => "10010000",
    1551 => "10010000",
    1552 => "10010000",
    1553 => "10010000",
    1554 => "10010000",
    1555 => "10010000",
    1556 => "10010000",
    1557 => "10010000",
    1558 => "10010000",
    1559 => "10010000",
    1560 => "10010000",
    1561 => "10010000",
    1562 => "10010000",
    1563 => "10010000",
    1564 => "10010000",
    1565 => "10010000",
    1566 => "10010000",
    1567 => "10010000",
    1568 => "10001111",
    1569 => "10001111",
    1570 => "10001111",
    1571 => "10001111",
    1572 => "10001111",
    1573 => "10001111",
    1574 => "10001111",
    1575 => "10001111",
    1576 => "10001111",
    1577 => "10001111",
    1578 => "10001111",
    1579 => "10001111",
    1580 => "10001111",
    1581 => "10001111",
    1582 => "10001111",
    1583 => "10001111",
    1584 => "10001111",
    1585 => "10001111",
    1586 => "10001111",
    1587 => "10001111",
    1588 => "10001111",
    1589 => "10001111",
    1590 => "10001111",
    1591 => "10001111",
    1592 => "10001111",
    1593 => "10001111",
    1594 => "10001111",
    1595 => "10001111",
    1596 => "10001111",
    1597 => "10001110",
    1598 => "10001110",
    1599 => "10001110",
    1600 => "10001110",
    1601 => "10001110",
    1602 => "10001110",
    1603 => "10001110",
    1604 => "10001110",
    1605 => "10001110",
    1606 => "10001110",
    1607 => "10001110",
    1608 => "10001110",
    1609 => "10001110",
    1610 => "10001110",
    1611 => "10001110",
    1612 => "10001110",
    1613 => "10001110",
    1614 => "10001110",
    1615 => "10001110",
    1616 => "10001110",
    1617 => "10001110",
    1618 => "10001110",
    1619 => "10001110",
    1620 => "10001110",
    1621 => "10001110",
    1622 => "10001110",
    1623 => "10001110",
    1624 => "10001110",
    1625 => "10001101",
    1626 => "10001101",
    1627 => "10001101",
    1628 => "10001101",
    1629 => "10001101",
    1630 => "10001101",
    1631 => "10001101",
    1632 => "10001101",
    1633 => "10001101",
    1634 => "10001101",
    1635 => "10001101",
    1636 => "10001101",
    1637 => "10001101",
    1638 => "10001101",
    1639 => "10001101",
    1640 => "10001101",
    1641 => "10001101",
    1642 => "10001101",
    1643 => "10001101",
    1644 => "10001101",
    1645 => "10001101",
    1646 => "10001101",
    1647 => "10001101",
    1648 => "10001101",
    1649 => "10001101",
    1650 => "10001101",
    1651 => "10001101",
    1652 => "10001101",
    1653 => "10001101",
    1654 => "10001100",
    1655 => "10001100",
    1656 => "10001100",
    1657 => "10001100",
    1658 => "10001100",
    1659 => "10001100",
    1660 => "10001100",
    1661 => "10001100",
    1662 => "10001100",
    1663 => "10001100",
    1664 => "10001100",
    1665 => "10001100",
    1666 => "10001100",
    1667 => "10001100",
    1668 => "10001100",
    1669 => "10001100",
    1670 => "10001100",
    1671 => "10001100",
    1672 => "10001100",
    1673 => "10001100",
    1674 => "10001100",
    1675 => "10001100",
    1676 => "10001100",
    1677 => "10001100",
    1678 => "10001100",
    1679 => "10001100",
    1680 => "10001100",
    1681 => "10001100",
    1682 => "10001011",
    1683 => "10001011",
    1684 => "10001011",
    1685 => "10001011",
    1686 => "10001011",
    1687 => "10001011",
    1688 => "10001011",
    1689 => "10001011",
    1690 => "10001011",
    1691 => "10001011",
    1692 => "10001011",
    1693 => "10001011",
    1694 => "10001011",
    1695 => "10001011",
    1696 => "10001011",
    1697 => "10001011",
    1698 => "10001011",
    1699 => "10001011",
    1700 => "10001011",
    1701 => "10001011",
    1702 => "10001011",
    1703 => "10001011",
    1704 => "10001011",
    1705 => "10001011",
    1706 => "10001011",
    1707 => "10001011",
    1708 => "10001011",
    1709 => "10001011",
    1710 => "10001011",
    1711 => "10001011",
    1712 => "10001010",
    1713 => "10001010",
    1714 => "10001010",
    1715 => "10001010",
    1716 => "10001010",
    1717 => "10001010",
    1718 => "10001010",
    1719 => "10001010",
    1720 => "10001010",
    1721 => "10001010",
    1722 => "10001010",
    1723 => "10001010",
    1724 => "10001010",
    1725 => "10001010",
    1726 => "10001010",
    1727 => "10001010",
    1728 => "10001010",
    1729 => "10001010",
    1730 => "10001010",
    1731 => "10001010",
    1732 => "10001010",
    1733 => "10001010",
    1734 => "10001010",
    1735 => "10001010",
    1736 => "10001010",
    1737 => "10001010",
    1738 => "10001010",
    1739 => "10001010",
    1740 => "10001010",
    1741 => "10001001",
    1742 => "10001001",
    1743 => "10001001",
    1744 => "10001001",
    1745 => "10001001",
    1746 => "10001001",
    1747 => "10001001",
    1748 => "10001001",
    1749 => "10001001",
    1750 => "10001001",
    1751 => "10001001",
    1752 => "10001001",
    1753 => "10001001",
    1754 => "10001001",
    1755 => "10001001",
    1756 => "10001001",
    1757 => "10001001",
    1758 => "10001001",
    1759 => "10001001",
    1760 => "10001001",
    1761 => "10001001",
    1762 => "10001001",
    1763 => "10001001",
    1764 => "10001001",
    1765 => "10001001",
    1766 => "10001001",
    1767 => "10001001",
    1768 => "10001001",
    1769 => "10001001",
    1770 => "10001001",
    1771 => "10001000",
    1772 => "10001000",
    1773 => "10001000",
    1774 => "10001000",
    1775 => "10001000",
    1776 => "10001000",
    1777 => "10001000",
    1778 => "10001000",
    1779 => "10001000",
    1780 => "10001000",
    1781 => "10001000",
    1782 => "10001000",
    1783 => "10001000",
    1784 => "10001000",
    1785 => "10001000",
    1786 => "10001000",
    1787 => "10001000",
    1788 => "10001000",
    1789 => "10001000",
    1790 => "10001000",
    1791 => "10001000",
    1792 => "10001000",
    1793 => "10001000",
    1794 => "10001000",
    1795 => "10001000",
    1796 => "10001000",
    1797 => "10001000",
    1798 => "10001000",
    1799 => "10001000",
    1800 => "10000111",
    1801 => "10000111",
    1802 => "10000111",
    1803 => "10000111",
    1804 => "10000111",
    1805 => "10000111",
    1806 => "10000111",
    1807 => "10000111",
    1808 => "10000111",
    1809 => "10000111",
    1810 => "10000111",
    1811 => "10000111",
    1812 => "10000111",
    1813 => "10000111",
    1814 => "10000111",
    1815 => "10000111",
    1816 => "10000111",
    1817 => "10000111",
    1818 => "10000111",
    1819 => "10000111",
    1820 => "10000111",
    1821 => "10000111",
    1822 => "10000111",
    1823 => "10000111",
    1824 => "10000111",
    1825 => "10000111",
    1826 => "10000111",
    1827 => "10000111",
    1828 => "10000111",
    1829 => "10000111",
    1830 => "10000111",
    1831 => "10000110",
    1832 => "10000110",
    1833 => "10000110",
    1834 => "10000110",
    1835 => "10000110",
    1836 => "10000110",
    1837 => "10000110",
    1838 => "10000110",
    1839 => "10000110",
    1840 => "10000110",
    1841 => "10000110",
    1842 => "10000110",
    1843 => "10000110",
    1844 => "10000110",
    1845 => "10000110",
    1846 => "10000110",
    1847 => "10000110",
    1848 => "10000110",
    1849 => "10000110",
    1850 => "10000110",
    1851 => "10000110",
    1852 => "10000110",
    1853 => "10000110",
    1854 => "10000110",
    1855 => "10000110",
    1856 => "10000110",
    1857 => "10000110",
    1858 => "10000110",
    1859 => "10000110",
    1860 => "10000110",
    1861 => "10000101",
    1862 => "10000101",
    1863 => "10000101",
    1864 => "10000101",
    1865 => "10000101",
    1866 => "10000101",
    1867 => "10000101",
    1868 => "10000101",
    1869 => "10000101",
    1870 => "10000101",
    1871 => "10000101",
    1872 => "10000101",
    1873 => "10000101",
    1874 => "10000101",
    1875 => "10000101",
    1876 => "10000101",
    1877 => "10000101",
    1878 => "10000101",
    1879 => "10000101",
    1880 => "10000101",
    1881 => "10000101",
    1882 => "10000101",
    1883 => "10000101",
    1884 => "10000101",
    1885 => "10000101",
    1886 => "10000101",
    1887 => "10000101",
    1888 => "10000101",
    1889 => "10000101",
    1890 => "10000101",
    1891 => "10000101",
    1892 => "10000100",
    1893 => "10000100",
    1894 => "10000100",
    1895 => "10000100",
    1896 => "10000100",
    1897 => "10000100",
    1898 => "10000100",
    1899 => "10000100",
    1900 => "10000100",
    1901 => "10000100",
    1902 => "10000100",
    1903 => "10000100",
    1904 => "10000100",
    1905 => "10000100",
    1906 => "10000100",
    1907 => "10000100",
    1908 => "10000100",
    1909 => "10000100",
    1910 => "10000100",
    1911 => "10000100",
    1912 => "10000100",
    1913 => "10000100",
    1914 => "10000100",
    1915 => "10000100",
    1916 => "10000100",
    1917 => "10000100",
    1918 => "10000100",
    1919 => "10000100",
    1920 => "10000100",
    1921 => "10000100",
    1922 => "10000011",
    1923 => "10000011",
    1924 => "10000011",
    1925 => "10000011",
    1926 => "10000011",
    1927 => "10000011",
    1928 => "10000011",
    1929 => "10000011",
    1930 => "10000011",
    1931 => "10000011",
    1932 => "10000011",
    1933 => "10000011",
    1934 => "10000011",
    1935 => "10000011",
    1936 => "10000011",
    1937 => "10000011",
    1938 => "10000011",
    1939 => "10000011",
    1940 => "10000011",
    1941 => "10000011",
    1942 => "10000011",
    1943 => "10000011",
    1944 => "10000011",
    1945 => "10000011",
    1946 => "10000011",
    1947 => "10000011",
    1948 => "10000011",
    1949 => "10000011",
    1950 => "10000011",
    1951 => "10000011",
    1952 => "10000011",
    1953 => "10000011",
    1954 => "10000010",
    1955 => "10000010",
    1956 => "10000010",
    1957 => "10000010",
    1958 => "10000010",
    1959 => "10000010",
    1960 => "10000010",
    1961 => "10000010",
    1962 => "10000010",
    1963 => "10000010",
    1964 => "10000010",
    1965 => "10000010",
    1966 => "10000010",
    1967 => "10000010",
    1968 => "10000010",
    1969 => "10000010",
    1970 => "10000010",
    1971 => "10000010",
    1972 => "10000010",
    1973 => "10000010",
    1974 => "10000010",
    1975 => "10000010",
    1976 => "10000010",
    1977 => "10000010",
    1978 => "10000010",
    1979 => "10000010",
    1980 => "10000010",
    1981 => "10000010",
    1982 => "10000010",
    1983 => "10000010",
    1984 => "10000010",
    1985 => "10000001",
    1986 => "10000001",
    1987 => "10000001",
    1988 => "10000001",
    1989 => "10000001",
    1990 => "10000001",
    1991 => "10000001",
    1992 => "10000001",
    1993 => "10000001",
    1994 => "10000001",
    1995 => "10000001",
    1996 => "10000001",
    1997 => "10000001",
    1998 => "10000001",
    1999 => "10000001",
    2000 => "10000001",
    2001 => "10000001",
    2002 => "10000001",
    2003 => "10000001",
    2004 => "10000001",
    2005 => "10000001",
    2006 => "10000001",
    2007 => "10000001",
    2008 => "10000001",
    2009 => "10000001",
    2010 => "10000001",
    2011 => "10000001",
    2012 => "10000001",
    2013 => "10000001",
    2014 => "10000001",
    2015 => "10000001",
    2016 => "10000001",
    2017 => "10000000",
    2018 => "10000000",
    2019 => "10000000",
    2020 => "10000000",
    2021 => "10000000",
    2022 => "10000000",
    2023 => "10000000",
    2024 => "10000000",
    2025 => "10000000",
    2026 => "10000000",
    2027 => "10000000",
    2028 => "10000000",
    2029 => "10000000",
    2030 => "10000000",
    2031 => "10000000",
    2032 => "10000000",
    2033 => "10000000",
    2034 => "10000000",
    2035 => "10000000",
    2036 => "10000000",
    2037 => "10000000",
    2038 => "10000000",
    2039 => "10000000",
    2040 => "10000000",
    2041 => "10000000",
    2042 => "10000000",
    2043 => "10000000",
    2044 => "10000000",
    2045 => "10000000",
    2046 => "10000000",
    2047 => "10000000",
    2048 => "01111111",
    2049 => "01111111",
    2050 => "01111111",
    2051 => "01111111",
    2052 => "01111111",
    2053 => "01111111",
    2054 => "01111111",
    2055 => "01111111",
    2056 => "01111111",
    2057 => "01111111",
    2058 => "01111111",
    2059 => "01111111",
    2060 => "01111111",
    2061 => "01111111",
    2062 => "01111111",
    2063 => "01111111",
    2064 => "01111111",
    2065 => "01111111",
    2066 => "01111111",
    2067 => "01111111",
    2068 => "01111111",
    2069 => "01111111",
    2070 => "01111111",
    2071 => "01111111",
    2072 => "01111111",
    2073 => "01111111",
    2074 => "01111111",
    2075 => "01111111",
    2076 => "01111111",
    2077 => "01111111",
    2078 => "01111111",
    2079 => "01111111",
    2080 => "01111111",
    2081 => "01111110",
    2082 => "01111110",
    2083 => "01111110",
    2084 => "01111110",
    2085 => "01111110",
    2086 => "01111110",
    2087 => "01111110",
    2088 => "01111110",
    2089 => "01111110",
    2090 => "01111110",
    2091 => "01111110",
    2092 => "01111110",
    2093 => "01111110",
    2094 => "01111110",
    2095 => "01111110",
    2096 => "01111110",
    2097 => "01111110",
    2098 => "01111110",
    2099 => "01111110",
    2100 => "01111110",
    2101 => "01111110",
    2102 => "01111110",
    2103 => "01111110",
    2104 => "01111110",
    2105 => "01111110",
    2106 => "01111110",
    2107 => "01111110",
    2108 => "01111110",
    2109 => "01111110",
    2110 => "01111110",
    2111 => "01111110",
    2112 => "01111110",
    2113 => "01111101",
    2114 => "01111101",
    2115 => "01111101",
    2116 => "01111101",
    2117 => "01111101",
    2118 => "01111101",
    2119 => "01111101",
    2120 => "01111101",
    2121 => "01111101",
    2122 => "01111101",
    2123 => "01111101",
    2124 => "01111101",
    2125 => "01111101",
    2126 => "01111101",
    2127 => "01111101",
    2128 => "01111101",
    2129 => "01111101",
    2130 => "01111101",
    2131 => "01111101",
    2132 => "01111101",
    2133 => "01111101",
    2134 => "01111101",
    2135 => "01111101",
    2136 => "01111101",
    2137 => "01111101",
    2138 => "01111101",
    2139 => "01111101",
    2140 => "01111101",
    2141 => "01111101",
    2142 => "01111101",
    2143 => "01111101",
    2144 => "01111101",
    2145 => "01111101",
    2146 => "01111100",
    2147 => "01111100",
    2148 => "01111100",
    2149 => "01111100",
    2150 => "01111100",
    2151 => "01111100",
    2152 => "01111100",
    2153 => "01111100",
    2154 => "01111100",
    2155 => "01111100",
    2156 => "01111100",
    2157 => "01111100",
    2158 => "01111100",
    2159 => "01111100",
    2160 => "01111100",
    2161 => "01111100",
    2162 => "01111100",
    2163 => "01111100",
    2164 => "01111100",
    2165 => "01111100",
    2166 => "01111100",
    2167 => "01111100",
    2168 => "01111100",
    2169 => "01111100",
    2170 => "01111100",
    2171 => "01111100",
    2172 => "01111100",
    2173 => "01111100",
    2174 => "01111100",
    2175 => "01111100",
    2176 => "01111100",
    2177 => "01111100",
    2178 => "01111011",
    2179 => "01111011",
    2180 => "01111011",
    2181 => "01111011",
    2182 => "01111011",
    2183 => "01111011",
    2184 => "01111011",
    2185 => "01111011",
    2186 => "01111011",
    2187 => "01111011",
    2188 => "01111011",
    2189 => "01111011",
    2190 => "01111011",
    2191 => "01111011",
    2192 => "01111011",
    2193 => "01111011",
    2194 => "01111011",
    2195 => "01111011",
    2196 => "01111011",
    2197 => "01111011",
    2198 => "01111011",
    2199 => "01111011",
    2200 => "01111011",
    2201 => "01111011",
    2202 => "01111011",
    2203 => "01111011",
    2204 => "01111011",
    2205 => "01111011",
    2206 => "01111011",
    2207 => "01111011",
    2208 => "01111011",
    2209 => "01111011",
    2210 => "01111011",
    2211 => "01111011",
    2212 => "01111010",
    2213 => "01111010",
    2214 => "01111010",
    2215 => "01111010",
    2216 => "01111010",
    2217 => "01111010",
    2218 => "01111010",
    2219 => "01111010",
    2220 => "01111010",
    2221 => "01111010",
    2222 => "01111010",
    2223 => "01111010",
    2224 => "01111010",
    2225 => "01111010",
    2226 => "01111010",
    2227 => "01111010",
    2228 => "01111010",
    2229 => "01111010",
    2230 => "01111010",
    2231 => "01111010",
    2232 => "01111010",
    2233 => "01111010",
    2234 => "01111010",
    2235 => "01111010",
    2236 => "01111010",
    2237 => "01111010",
    2238 => "01111010",
    2239 => "01111010",
    2240 => "01111010",
    2241 => "01111010",
    2242 => "01111010",
    2243 => "01111010",
    2244 => "01111010",
    2245 => "01111001",
    2246 => "01111001",
    2247 => "01111001",
    2248 => "01111001",
    2249 => "01111001",
    2250 => "01111001",
    2251 => "01111001",
    2252 => "01111001",
    2253 => "01111001",
    2254 => "01111001",
    2255 => "01111001",
    2256 => "01111001",
    2257 => "01111001",
    2258 => "01111001",
    2259 => "01111001",
    2260 => "01111001",
    2261 => "01111001",
    2262 => "01111001",
    2263 => "01111001",
    2264 => "01111001",
    2265 => "01111001",
    2266 => "01111001",
    2267 => "01111001",
    2268 => "01111001",
    2269 => "01111001",
    2270 => "01111001",
    2271 => "01111001",
    2272 => "01111001",
    2273 => "01111001",
    2274 => "01111001",
    2275 => "01111001",
    2276 => "01111001",
    2277 => "01111001",
    2278 => "01111001",
    2279 => "01111000",
    2280 => "01111000",
    2281 => "01111000",
    2282 => "01111000",
    2283 => "01111000",
    2284 => "01111000",
    2285 => "01111000",
    2286 => "01111000",
    2287 => "01111000",
    2288 => "01111000",
    2289 => "01111000",
    2290 => "01111000",
    2291 => "01111000",
    2292 => "01111000",
    2293 => "01111000",
    2294 => "01111000",
    2295 => "01111000",
    2296 => "01111000",
    2297 => "01111000",
    2298 => "01111000",
    2299 => "01111000",
    2300 => "01111000",
    2301 => "01111000",
    2302 => "01111000",
    2303 => "01111000",
    2304 => "01111000",
    2305 => "01111000",
    2306 => "01111000",
    2307 => "01111000",
    2308 => "01111000",
    2309 => "01111000",
    2310 => "01111000",
    2311 => "01111000",
    2312 => "01110111",
    2313 => "01110111",
    2314 => "01110111",
    2315 => "01110111",
    2316 => "01110111",
    2317 => "01110111",
    2318 => "01110111",
    2319 => "01110111",
    2320 => "01110111",
    2321 => "01110111",
    2322 => "01110111",
    2323 => "01110111",
    2324 => "01110111",
    2325 => "01110111",
    2326 => "01110111",
    2327 => "01110111",
    2328 => "01110111",
    2329 => "01110111",
    2330 => "01110111",
    2331 => "01110111",
    2332 => "01110111",
    2333 => "01110111",
    2334 => "01110111",
    2335 => "01110111",
    2336 => "01110111",
    2337 => "01110111",
    2338 => "01110111",
    2339 => "01110111",
    2340 => "01110111",
    2341 => "01110111",
    2342 => "01110111",
    2343 => "01110111",
    2344 => "01110111",
    2345 => "01110111",
    2346 => "01110111",
    2347 => "01110110",
    2348 => "01110110",
    2349 => "01110110",
    2350 => "01110110",
    2351 => "01110110",
    2352 => "01110110",
    2353 => "01110110",
    2354 => "01110110",
    2355 => "01110110",
    2356 => "01110110",
    2357 => "01110110",
    2358 => "01110110",
    2359 => "01110110",
    2360 => "01110110",
    2361 => "01110110",
    2362 => "01110110",
    2363 => "01110110",
    2364 => "01110110",
    2365 => "01110110",
    2366 => "01110110",
    2367 => "01110110",
    2368 => "01110110",
    2369 => "01110110",
    2370 => "01110110",
    2371 => "01110110",
    2372 => "01110110",
    2373 => "01110110",
    2374 => "01110110",
    2375 => "01110110",
    2376 => "01110110",
    2377 => "01110110",
    2378 => "01110110",
    2379 => "01110110",
    2380 => "01110110",
    2381 => "01110101",
    2382 => "01110101",
    2383 => "01110101",
    2384 => "01110101",
    2385 => "01110101",
    2386 => "01110101",
    2387 => "01110101",
    2388 => "01110101",
    2389 => "01110101",
    2390 => "01110101",
    2391 => "01110101",
    2392 => "01110101",
    2393 => "01110101",
    2394 => "01110101",
    2395 => "01110101",
    2396 => "01110101",
    2397 => "01110101",
    2398 => "01110101",
    2399 => "01110101",
    2400 => "01110101",
    2401 => "01110101",
    2402 => "01110101",
    2403 => "01110101",
    2404 => "01110101",
    2405 => "01110101",
    2406 => "01110101",
    2407 => "01110101",
    2408 => "01110101",
    2409 => "01110101",
    2410 => "01110101",
    2411 => "01110101",
    2412 => "01110101",
    2413 => "01110101",
    2414 => "01110101",
    2415 => "01110101",
    2416 => "01110100",
    2417 => "01110100",
    2418 => "01110100",
    2419 => "01110100",
    2420 => "01110100",
    2421 => "01110100",
    2422 => "01110100",
    2423 => "01110100",
    2424 => "01110100",
    2425 => "01110100",
    2426 => "01110100",
    2427 => "01110100",
    2428 => "01110100",
    2429 => "01110100",
    2430 => "01110100",
    2431 => "01110100",
    2432 => "01110100",
    2433 => "01110100",
    2434 => "01110100",
    2435 => "01110100",
    2436 => "01110100",
    2437 => "01110100",
    2438 => "01110100",
    2439 => "01110100",
    2440 => "01110100",
    2441 => "01110100",
    2442 => "01110100",
    2443 => "01110100",
    2444 => "01110100",
    2445 => "01110100",
    2446 => "01110100",
    2447 => "01110100",
    2448 => "01110100",
    2449 => "01110100",
    2450 => "01110011",
    2451 => "01110011",
    2452 => "01110011",
    2453 => "01110011",
    2454 => "01110011",
    2455 => "01110011",
    2456 => "01110011",
    2457 => "01110011",
    2458 => "01110011",
    2459 => "01110011",
    2460 => "01110011",
    2461 => "01110011",
    2462 => "01110011",
    2463 => "01110011",
    2464 => "01110011",
    2465 => "01110011",
    2466 => "01110011",
    2467 => "01110011",
    2468 => "01110011",
    2469 => "01110011",
    2470 => "01110011",
    2471 => "01110011",
    2472 => "01110011",
    2473 => "01110011",
    2474 => "01110011",
    2475 => "01110011",
    2476 => "01110011",
    2477 => "01110011",
    2478 => "01110011",
    2479 => "01110011",
    2480 => "01110011",
    2481 => "01110011",
    2482 => "01110011",
    2483 => "01110011",
    2484 => "01110011",
    2485 => "01110011",
    2486 => "01110010",
    2487 => "01110010",
    2488 => "01110010",
    2489 => "01110010",
    2490 => "01110010",
    2491 => "01110010",
    2492 => "01110010",
    2493 => "01110010",
    2494 => "01110010",
    2495 => "01110010",
    2496 => "01110010",
    2497 => "01110010",
    2498 => "01110010",
    2499 => "01110010",
    2500 => "01110010",
    2501 => "01110010",
    2502 => "01110010",
    2503 => "01110010",
    2504 => "01110010",
    2505 => "01110010",
    2506 => "01110010",
    2507 => "01110010",
    2508 => "01110010",
    2509 => "01110010",
    2510 => "01110010",
    2511 => "01110010",
    2512 => "01110010",
    2513 => "01110010",
    2514 => "01110010",
    2515 => "01110010",
    2516 => "01110010",
    2517 => "01110010",
    2518 => "01110010",
    2519 => "01110010",
    2520 => "01110010",
    2521 => "01110001",
    2522 => "01110001",
    2523 => "01110001",
    2524 => "01110001",
    2525 => "01110001",
    2526 => "01110001",
    2527 => "01110001",
    2528 => "01110001",
    2529 => "01110001",
    2530 => "01110001",
    2531 => "01110001",
    2532 => "01110001",
    2533 => "01110001",
    2534 => "01110001",
    2535 => "01110001",
    2536 => "01110001",
    2537 => "01110001",
    2538 => "01110001",
    2539 => "01110001",
    2540 => "01110001",
    2541 => "01110001",
    2542 => "01110001",
    2543 => "01110001",
    2544 => "01110001",
    2545 => "01110001",
    2546 => "01110001",
    2547 => "01110001",
    2548 => "01110001",
    2549 => "01110001",
    2550 => "01110001",
    2551 => "01110001",
    2552 => "01110001",
    2553 => "01110001",
    2554 => "01110001",
    2555 => "01110001",
    2556 => "01110001",
    2557 => "01110000",
    2558 => "01110000",
    2559 => "01110000",
    2560 => "01110000",
    2561 => "01110000",
    2562 => "01110000",
    2563 => "01110000",
    2564 => "01110000",
    2565 => "01110000",
    2566 => "01110000",
    2567 => "01110000",
    2568 => "01110000",
    2569 => "01110000",
    2570 => "01110000",
    2571 => "01110000",
    2572 => "01110000",
    2573 => "01110000",
    2574 => "01110000",
    2575 => "01110000",
    2576 => "01110000",
    2577 => "01110000",
    2578 => "01110000",
    2579 => "01110000",
    2580 => "01110000",
    2581 => "01110000",
    2582 => "01110000",
    2583 => "01110000",
    2584 => "01110000",
    2585 => "01110000",
    2586 => "01110000",
    2587 => "01110000",
    2588 => "01110000",
    2589 => "01110000",
    2590 => "01110000",
    2591 => "01110000",
    2592 => "01101111",
    2593 => "01101111",
    2594 => "01101111",
    2595 => "01101111",
    2596 => "01101111",
    2597 => "01101111",
    2598 => "01101111",
    2599 => "01101111",
    2600 => "01101111",
    2601 => "01101111",
    2602 => "01101111",
    2603 => "01101111",
    2604 => "01101111",
    2605 => "01101111",
    2606 => "01101111",
    2607 => "01101111",
    2608 => "01101111",
    2609 => "01101111",
    2610 => "01101111",
    2611 => "01101111",
    2612 => "01101111",
    2613 => "01101111",
    2614 => "01101111",
    2615 => "01101111",
    2616 => "01101111",
    2617 => "01101111",
    2618 => "01101111",
    2619 => "01101111",
    2620 => "01101111",
    2621 => "01101111",
    2622 => "01101111",
    2623 => "01101111",
    2624 => "01101111",
    2625 => "01101111",
    2626 => "01101111",
    2627 => "01101111",
    2628 => "01101111",
    2629 => "01101110",
    2630 => "01101110",
    2631 => "01101110",
    2632 => "01101110",
    2633 => "01101110",
    2634 => "01101110",
    2635 => "01101110",
    2636 => "01101110",
    2637 => "01101110",
    2638 => "01101110",
    2639 => "01101110",
    2640 => "01101110",
    2641 => "01101110",
    2642 => "01101110",
    2643 => "01101110",
    2644 => "01101110",
    2645 => "01101110",
    2646 => "01101110",
    2647 => "01101110",
    2648 => "01101110",
    2649 => "01101110",
    2650 => "01101110",
    2651 => "01101110",
    2652 => "01101110",
    2653 => "01101110",
    2654 => "01101110",
    2655 => "01101110",
    2656 => "01101110",
    2657 => "01101110",
    2658 => "01101110",
    2659 => "01101110",
    2660 => "01101110",
    2661 => "01101110",
    2662 => "01101110",
    2663 => "01101110",
    2664 => "01101110",
    2665 => "01101101",
    2666 => "01101101",
    2667 => "01101101",
    2668 => "01101101",
    2669 => "01101101",
    2670 => "01101101",
    2671 => "01101101",
    2672 => "01101101",
    2673 => "01101101",
    2674 => "01101101",
    2675 => "01101101",
    2676 => "01101101",
    2677 => "01101101",
    2678 => "01101101",
    2679 => "01101101",
    2680 => "01101101",
    2681 => "01101101",
    2682 => "01101101",
    2683 => "01101101",
    2684 => "01101101",
    2685 => "01101101",
    2686 => "01101101",
    2687 => "01101101",
    2688 => "01101101",
    2689 => "01101101",
    2690 => "01101101",
    2691 => "01101101",
    2692 => "01101101",
    2693 => "01101101",
    2694 => "01101101",
    2695 => "01101101",
    2696 => "01101101",
    2697 => "01101101",
    2698 => "01101101",
    2699 => "01101101",
    2700 => "01101101",
    2701 => "01101101",
    2702 => "01101100",
    2703 => "01101100",
    2704 => "01101100",
    2705 => "01101100",
    2706 => "01101100",
    2707 => "01101100",
    2708 => "01101100",
    2709 => "01101100",
    2710 => "01101100",
    2711 => "01101100",
    2712 => "01101100",
    2713 => "01101100",
    2714 => "01101100",
    2715 => "01101100",
    2716 => "01101100",
    2717 => "01101100",
    2718 => "01101100",
    2719 => "01101100",
    2720 => "01101100",
    2721 => "01101100",
    2722 => "01101100",
    2723 => "01101100",
    2724 => "01101100",
    2725 => "01101100",
    2726 => "01101100",
    2727 => "01101100",
    2728 => "01101100",
    2729 => "01101100",
    2730 => "01101100",
    2731 => "01101100",
    2732 => "01101100",
    2733 => "01101100",
    2734 => "01101100",
    2735 => "01101100",
    2736 => "01101100",
    2737 => "01101100",
    2738 => "01101011",
    2739 => "01101011",
    2740 => "01101011",
    2741 => "01101011",
    2742 => "01101011",
    2743 => "01101011",
    2744 => "01101011",
    2745 => "01101011",
    2746 => "01101011",
    2747 => "01101011",
    2748 => "01101011",
    2749 => "01101011",
    2750 => "01101011",
    2751 => "01101011",
    2752 => "01101011",
    2753 => "01101011",
    2754 => "01101011",
    2755 => "01101011",
    2756 => "01101011",
    2757 => "01101011",
    2758 => "01101011",
    2759 => "01101011",
    2760 => "01101011",
    2761 => "01101011",
    2762 => "01101011",
    2763 => "01101011",
    2764 => "01101011",
    2765 => "01101011",
    2766 => "01101011",
    2767 => "01101011",
    2768 => "01101011",
    2769 => "01101011",
    2770 => "01101011",
    2771 => "01101011",
    2772 => "01101011",
    2773 => "01101011",
    2774 => "01101011",
    2775 => "01101011",
    2776 => "01101010",
    2777 => "01101010",
    2778 => "01101010",
    2779 => "01101010",
    2780 => "01101010",
    2781 => "01101010",
    2782 => "01101010",
    2783 => "01101010",
    2784 => "01101010",
    2785 => "01101010",
    2786 => "01101010",
    2787 => "01101010",
    2788 => "01101010",
    2789 => "01101010",
    2790 => "01101010",
    2791 => "01101010",
    2792 => "01101010",
    2793 => "01101010",
    2794 => "01101010",
    2795 => "01101010",
    2796 => "01101010",
    2797 => "01101010",
    2798 => "01101010",
    2799 => "01101010",
    2800 => "01101010",
    2801 => "01101010",
    2802 => "01101010",
    2803 => "01101010",
    2804 => "01101010",
    2805 => "01101010",
    2806 => "01101010",
    2807 => "01101010",
    2808 => "01101010",
    2809 => "01101010",
    2810 => "01101010",
    2811 => "01101010",
    2812 => "01101010",
    2813 => "01101001",
    2814 => "01101001",
    2815 => "01101001",
    2816 => "01101001",
    2817 => "01101001",
    2818 => "01101001",
    2819 => "01101001",
    2820 => "01101001",
    2821 => "01101001",
    2822 => "01101001",
    2823 => "01101001",
    2824 => "01101001",
    2825 => "01101001",
    2826 => "01101001",
    2827 => "01101001",
    2828 => "01101001",
    2829 => "01101001",
    2830 => "01101001",
    2831 => "01101001",
    2832 => "01101001",
    2833 => "01101001",
    2834 => "01101001",
    2835 => "01101001",
    2836 => "01101001",
    2837 => "01101001",
    2838 => "01101001",
    2839 => "01101001",
    2840 => "01101001",
    2841 => "01101001",
    2842 => "01101001",
    2843 => "01101001",
    2844 => "01101001",
    2845 => "01101001",
    2846 => "01101001",
    2847 => "01101001",
    2848 => "01101001",
    2849 => "01101001",
    2850 => "01101001",
    2851 => "01101000",
    2852 => "01101000",
    2853 => "01101000",
    2854 => "01101000",
    2855 => "01101000",
    2856 => "01101000",
    2857 => "01101000",
    2858 => "01101000",
    2859 => "01101000",
    2860 => "01101000",
    2861 => "01101000",
    2862 => "01101000",
    2863 => "01101000",
    2864 => "01101000",
    2865 => "01101000",
    2866 => "01101000",
    2867 => "01101000",
    2868 => "01101000",
    2869 => "01101000",
    2870 => "01101000",
    2871 => "01101000",
    2872 => "01101000",
    2873 => "01101000",
    2874 => "01101000",
    2875 => "01101000",
    2876 => "01101000",
    2877 => "01101000",
    2878 => "01101000",
    2879 => "01101000",
    2880 => "01101000",
    2881 => "01101000",
    2882 => "01101000",
    2883 => "01101000",
    2884 => "01101000",
    2885 => "01101000",
    2886 => "01101000",
    2887 => "01101000",
    2888 => "01100111",
    2889 => "01100111",
    2890 => "01100111",
    2891 => "01100111",
    2892 => "01100111",
    2893 => "01100111",
    2894 => "01100111",
    2895 => "01100111",
    2896 => "01100111",
    2897 => "01100111",
    2898 => "01100111",
    2899 => "01100111",
    2900 => "01100111",
    2901 => "01100111",
    2902 => "01100111",
    2903 => "01100111",
    2904 => "01100111",
    2905 => "01100111",
    2906 => "01100111",
    2907 => "01100111",
    2908 => "01100111",
    2909 => "01100111",
    2910 => "01100111",
    2911 => "01100111",
    2912 => "01100111",
    2913 => "01100111",
    2914 => "01100111",
    2915 => "01100111",
    2916 => "01100111",
    2917 => "01100111",
    2918 => "01100111",
    2919 => "01100111",
    2920 => "01100111",
    2921 => "01100111",
    2922 => "01100111",
    2923 => "01100111",
    2924 => "01100111",
    2925 => "01100111",
    2926 => "01100111",
    2927 => "01100110",
    2928 => "01100110",
    2929 => "01100110",
    2930 => "01100110",
    2931 => "01100110",
    2932 => "01100110",
    2933 => "01100110",
    2934 => "01100110",
    2935 => "01100110",
    2936 => "01100110",
    2937 => "01100110",
    2938 => "01100110",
    2939 => "01100110",
    2940 => "01100110",
    2941 => "01100110",
    2942 => "01100110",
    2943 => "01100110",
    2944 => "01100110",
    2945 => "01100110",
    2946 => "01100110",
    2947 => "01100110",
    2948 => "01100110",
    2949 => "01100110",
    2950 => "01100110",
    2951 => "01100110",
    2952 => "01100110",
    2953 => "01100110",
    2954 => "01100110",
    2955 => "01100110",
    2956 => "01100110",
    2957 => "01100110",
    2958 => "01100110",
    2959 => "01100110",
    2960 => "01100110",
    2961 => "01100110",
    2962 => "01100110",
    2963 => "01100110",
    2964 => "01100110",
    2965 => "01100101",
    2966 => "01100101",
    2967 => "01100101",
    2968 => "01100101",
    2969 => "01100101",
    2970 => "01100101",
    2971 => "01100101",
    2972 => "01100101",
    2973 => "01100101",
    2974 => "01100101",
    2975 => "01100101",
    2976 => "01100101",
    2977 => "01100101",
    2978 => "01100101",
    2979 => "01100101",
    2980 => "01100101",
    2981 => "01100101",
    2982 => "01100101",
    2983 => "01100101",
    2984 => "01100101",
    2985 => "01100101",
    2986 => "01100101",
    2987 => "01100101",
    2988 => "01100101",
    2989 => "01100101",
    2990 => "01100101",
    2991 => "01100101",
    2992 => "01100101",
    2993 => "01100101",
    2994 => "01100101",
    2995 => "01100101",
    2996 => "01100101",
    2997 => "01100101",
    2998 => "01100101",
    2999 => "01100101",
    3000 => "01100101",
    3001 => "01100101",
    3002 => "01100101",
    3003 => "01100101",
    3004 => "01100100",
    3005 => "01100100",
    3006 => "01100100",
    3007 => "01100100",
    3008 => "01100100",
    3009 => "01100100",
    3010 => "01100100",
    3011 => "01100100",
    3012 => "01100100",
    3013 => "01100100",
    3014 => "01100100",
    3015 => "01100100",
    3016 => "01100100",
    3017 => "01100100",
    3018 => "01100100",
    3019 => "01100100",
    3020 => "01100100",
    3021 => "01100100",
    3022 => "01100100",
    3023 => "01100100",
    3024 => "01100100",
    3025 => "01100100",
    3026 => "01100100",
    3027 => "01100100",
    3028 => "01100100",
    3029 => "01100100",
    3030 => "01100100",
    3031 => "01100100",
    3032 => "01100100",
    3033 => "01100100",
    3034 => "01100100",
    3035 => "01100100",
    3036 => "01100100",
    3037 => "01100100",
    3038 => "01100100",
    3039 => "01100100",
    3040 => "01100100",
    3041 => "01100100",
    3042 => "01100011",
    3043 => "01100011",
    3044 => "01100011",
    3045 => "01100011",
    3046 => "01100011",
    3047 => "01100011",
    3048 => "01100011",
    3049 => "01100011",
    3050 => "01100011",
    3051 => "01100011",
    3052 => "01100011",
    3053 => "01100011",
    3054 => "01100011",
    3055 => "01100011",
    3056 => "01100011",
    3057 => "01100011",
    3058 => "01100011",
    3059 => "01100011",
    3060 => "01100011",
    3061 => "01100011",
    3062 => "01100011",
    3063 => "01100011",
    3064 => "01100011",
    3065 => "01100011",
    3066 => "01100011",
    3067 => "01100011",
    3068 => "01100011",
    3069 => "01100011",
    3070 => "01100011",
    3071 => "01100011",
    3072 => "01100011",
    3073 => "01100011",
    3074 => "01100011",
    3075 => "01100011",
    3076 => "01100011",
    3077 => "01100011",
    3078 => "01100011",
    3079 => "01100011",
    3080 => "01100011",
    3081 => "01100011",
    3082 => "01100010",
    3083 => "01100010",
    3084 => "01100010",
    3085 => "01100010",
    3086 => "01100010",
    3087 => "01100010",
    3088 => "01100010",
    3089 => "01100010",
    3090 => "01100010",
    3091 => "01100010",
    3092 => "01100010",
    3093 => "01100010",
    3094 => "01100010",
    3095 => "01100010",
    3096 => "01100010",
    3097 => "01100010",
    3098 => "01100010",
    3099 => "01100010",
    3100 => "01100010",
    3101 => "01100010",
    3102 => "01100010",
    3103 => "01100010",
    3104 => "01100010",
    3105 => "01100010",
    3106 => "01100010",
    3107 => "01100010",
    3108 => "01100010",
    3109 => "01100010",
    3110 => "01100010",
    3111 => "01100010",
    3112 => "01100010",
    3113 => "01100010",
    3114 => "01100010",
    3115 => "01100010",
    3116 => "01100010",
    3117 => "01100010",
    3118 => "01100010",
    3119 => "01100010",
    3120 => "01100010",
    3121 => "01100001",
    3122 => "01100001",
    3123 => "01100001",
    3124 => "01100001",
    3125 => "01100001",
    3126 => "01100001",
    3127 => "01100001",
    3128 => "01100001",
    3129 => "01100001",
    3130 => "01100001",
    3131 => "01100001",
    3132 => "01100001",
    3133 => "01100001",
    3134 => "01100001",
    3135 => "01100001",
    3136 => "01100001",
    3137 => "01100001",
    3138 => "01100001",
    3139 => "01100001",
    3140 => "01100001",
    3141 => "01100001",
    3142 => "01100001",
    3143 => "01100001",
    3144 => "01100001",
    3145 => "01100001",
    3146 => "01100001",
    3147 => "01100001",
    3148 => "01100001",
    3149 => "01100001",
    3150 => "01100001",
    3151 => "01100001",
    3152 => "01100001",
    3153 => "01100001",
    3154 => "01100001",
    3155 => "01100001",
    3156 => "01100001",
    3157 => "01100001",
    3158 => "01100001",
    3159 => "01100001",
    3160 => "01100001",
    3161 => "01100000",
    3162 => "01100000",
    3163 => "01100000",
    3164 => "01100000",
    3165 => "01100000",
    3166 => "01100000",
    3167 => "01100000",
    3168 => "01100000",
    3169 => "01100000",
    3170 => "01100000",
    3171 => "01100000",
    3172 => "01100000",
    3173 => "01100000",
    3174 => "01100000",
    3175 => "01100000",
    3176 => "01100000",
    3177 => "01100000",
    3178 => "01100000",
    3179 => "01100000",
    3180 => "01100000",
    3181 => "01100000",
    3182 => "01100000",
    3183 => "01100000",
    3184 => "01100000",
    3185 => "01100000",
    3186 => "01100000",
    3187 => "01100000",
    3188 => "01100000",
    3189 => "01100000",
    3190 => "01100000",
    3191 => "01100000",
    3192 => "01100000",
    3193 => "01100000",
    3194 => "01100000",
    3195 => "01100000",
    3196 => "01100000",
    3197 => "01100000",
    3198 => "01100000",
    3199 => "01100000",
    3200 => "01011111",
    3201 => "01011111",
    3202 => "01011111",
    3203 => "01011111",
    3204 => "01011111",
    3205 => "01011111",
    3206 => "01011111",
    3207 => "01011111",
    3208 => "01011111",
    3209 => "01011111",
    3210 => "01011111",
    3211 => "01011111",
    3212 => "01011111",
    3213 => "01011111",
    3214 => "01011111",
    3215 => "01011111",
    3216 => "01011111",
    3217 => "01011111",
    3218 => "01011111",
    3219 => "01011111",
    3220 => "01011111",
    3221 => "01011111",
    3222 => "01011111",
    3223 => "01011111",
    3224 => "01011111",
    3225 => "01011111",
    3226 => "01011111",
    3227 => "01011111",
    3228 => "01011111",
    3229 => "01011111",
    3230 => "01011111",
    3231 => "01011111",
    3232 => "01011111",
    3233 => "01011111",
    3234 => "01011111",
    3235 => "01011111",
    3236 => "01011111",
    3237 => "01011111",
    3238 => "01011111",
    3239 => "01011111",
    3240 => "01011111",
    3241 => "01011110",
    3242 => "01011110",
    3243 => "01011110",
    3244 => "01011110",
    3245 => "01011110",
    3246 => "01011110",
    3247 => "01011110",
    3248 => "01011110",
    3249 => "01011110",
    3250 => "01011110",
    3251 => "01011110",
    3252 => "01011110",
    3253 => "01011110",
    3254 => "01011110",
    3255 => "01011110",
    3256 => "01011110",
    3257 => "01011110",
    3258 => "01011110",
    3259 => "01011110",
    3260 => "01011110",
    3261 => "01011110",
    3262 => "01011110",
    3263 => "01011110",
    3264 => "01011110",
    3265 => "01011110",
    3266 => "01011110",
    3267 => "01011110",
    3268 => "01011110",
    3269 => "01011110",
    3270 => "01011110",
    3271 => "01011110",
    3272 => "01011110",
    3273 => "01011110",
    3274 => "01011110",
    3275 => "01011110",
    3276 => "01011110",
    3277 => "01011110",
    3278 => "01011110",
    3279 => "01011110",
    3280 => "01011110",
    3281 => "01011101",
    3282 => "01011101",
    3283 => "01011101",
    3284 => "01011101",
    3285 => "01011101",
    3286 => "01011101",
    3287 => "01011101",
    3288 => "01011101",
    3289 => "01011101",
    3290 => "01011101",
    3291 => "01011101",
    3292 => "01011101",
    3293 => "01011101",
    3294 => "01011101",
    3295 => "01011101",
    3296 => "01011101",
    3297 => "01011101",
    3298 => "01011101",
    3299 => "01011101",
    3300 => "01011101",
    3301 => "01011101",
    3302 => "01011101",
    3303 => "01011101",
    3304 => "01011101",
    3305 => "01011101",
    3306 => "01011101",
    3307 => "01011101",
    3308 => "01011101",
    3309 => "01011101",
    3310 => "01011101",
    3311 => "01011101",
    3312 => "01011101",
    3313 => "01011101",
    3314 => "01011101",
    3315 => "01011101",
    3316 => "01011101",
    3317 => "01011101",
    3318 => "01011101",
    3319 => "01011101",
    3320 => "01011101",
    3321 => "01011101",
    3322 => "01011100",
    3323 => "01011100",
    3324 => "01011100",
    3325 => "01011100",
    3326 => "01011100",
    3327 => "01011100",
    3328 => "01011100",
    3329 => "01011100",
    3330 => "01011100",
    3331 => "01011100",
    3332 => "01011100",
    3333 => "01011100",
    3334 => "01011100",
    3335 => "01011100",
    3336 => "01011100",
    3337 => "01011100",
    3338 => "01011100",
    3339 => "01011100",
    3340 => "01011100",
    3341 => "01011100",
    3342 => "01011100",
    3343 => "01011100",
    3344 => "01011100",
    3345 => "01011100",
    3346 => "01011100",
    3347 => "01011100",
    3348 => "01011100",
    3349 => "01011100",
    3350 => "01011100",
    3351 => "01011100",
    3352 => "01011100",
    3353 => "01011100",
    3354 => "01011100",
    3355 => "01011100",
    3356 => "01011100",
    3357 => "01011100",
    3358 => "01011100",
    3359 => "01011100",
    3360 => "01011100",
    3361 => "01011100",
    3362 => "01011011",
    3363 => "01011011",
    3364 => "01011011",
    3365 => "01011011",
    3366 => "01011011",
    3367 => "01011011",
    3368 => "01011011",
    3369 => "01011011",
    3370 => "01011011",
    3371 => "01011011",
    3372 => "01011011",
    3373 => "01011011",
    3374 => "01011011",
    3375 => "01011011",
    3376 => "01011011",
    3377 => "01011011",
    3378 => "01011011",
    3379 => "01011011",
    3380 => "01011011",
    3381 => "01011011",
    3382 => "01011011",
    3383 => "01011011",
    3384 => "01011011",
    3385 => "01011011",
    3386 => "01011011",
    3387 => "01011011",
    3388 => "01011011",
    3389 => "01011011",
    3390 => "01011011",
    3391 => "01011011",
    3392 => "01011011",
    3393 => "01011011",
    3394 => "01011011",
    3395 => "01011011",
    3396 => "01011011",
    3397 => "01011011",
    3398 => "01011011",
    3399 => "01011011",
    3400 => "01011011",
    3401 => "01011011",
    3402 => "01011011",
    3403 => "01011011",
    3404 => "01011010",
    3405 => "01011010",
    3406 => "01011010",
    3407 => "01011010",
    3408 => "01011010",
    3409 => "01011010",
    3410 => "01011010",
    3411 => "01011010",
    3412 => "01011010",
    3413 => "01011010",
    3414 => "01011010",
    3415 => "01011010",
    3416 => "01011010",
    3417 => "01011010",
    3418 => "01011010",
    3419 => "01011010",
    3420 => "01011010",
    3421 => "01011010",
    3422 => "01011010",
    3423 => "01011010",
    3424 => "01011010",
    3425 => "01011010",
    3426 => "01011010",
    3427 => "01011010",
    3428 => "01011010",
    3429 => "01011010",
    3430 => "01011010",
    3431 => "01011010",
    3432 => "01011010",
    3433 => "01011010",
    3434 => "01011010",
    3435 => "01011010",
    3436 => "01011010",
    3437 => "01011010",
    3438 => "01011010",
    3439 => "01011010",
    3440 => "01011010",
    3441 => "01011010",
    3442 => "01011010",
    3443 => "01011010",
    3444 => "01011010",
    3445 => "01011001",
    3446 => "01011001",
    3447 => "01011001",
    3448 => "01011001",
    3449 => "01011001",
    3450 => "01011001",
    3451 => "01011001",
    3452 => "01011001",
    3453 => "01011001",
    3454 => "01011001",
    3455 => "01011001",
    3456 => "01011001",
    3457 => "01011001",
    3458 => "01011001",
    3459 => "01011001",
    3460 => "01011001",
    3461 => "01011001",
    3462 => "01011001",
    3463 => "01011001",
    3464 => "01011001",
    3465 => "01011001",
    3466 => "01011001",
    3467 => "01011001",
    3468 => "01011001",
    3469 => "01011001",
    3470 => "01011001",
    3471 => "01011001",
    3472 => "01011001",
    3473 => "01011001",
    3474 => "01011001",
    3475 => "01011001",
    3476 => "01011001",
    3477 => "01011001",
    3478 => "01011001",
    3479 => "01011001",
    3480 => "01011001",
    3481 => "01011001",
    3482 => "01011001",
    3483 => "01011001",
    3484 => "01011001",
    3485 => "01011001",
    3486 => "01011001",
    3487 => "01011000",
    3488 => "01011000",
    3489 => "01011000",
    3490 => "01011000",
    3491 => "01011000",
    3492 => "01011000",
    3493 => "01011000",
    3494 => "01011000",
    3495 => "01011000",
    3496 => "01011000",
    3497 => "01011000",
    3498 => "01011000",
    3499 => "01011000",
    3500 => "01011000",
    3501 => "01011000",
    3502 => "01011000",
    3503 => "01011000",
    3504 => "01011000",
    3505 => "01011000",
    3506 => "01011000",
    3507 => "01011000",
    3508 => "01011000",
    3509 => "01011000",
    3510 => "01011000",
    3511 => "01011000",
    3512 => "01011000",
    3513 => "01011000",
    3514 => "01011000",
    3515 => "01011000",
    3516 => "01011000",
    3517 => "01011000",
    3518 => "01011000",
    3519 => "01011000",
    3520 => "01011000",
    3521 => "01011000",
    3522 => "01011000",
    3523 => "01011000",
    3524 => "01011000",
    3525 => "01011000",
    3526 => "01011000",
    3527 => "01011000",
    3528 => "01010111",
    3529 => "01010111",
    3530 => "01010111",
    3531 => "01010111",
    3532 => "01010111",
    3533 => "01010111",
    3534 => "01010111",
    3535 => "01010111",
    3536 => "01010111",
    3537 => "01010111",
    3538 => "01010111",
    3539 => "01010111",
    3540 => "01010111",
    3541 => "01010111",
    3542 => "01010111",
    3543 => "01010111",
    3544 => "01010111",
    3545 => "01010111",
    3546 => "01010111",
    3547 => "01010111",
    3548 => "01010111",
    3549 => "01010111",
    3550 => "01010111",
    3551 => "01010111",
    3552 => "01010111",
    3553 => "01010111",
    3554 => "01010111",
    3555 => "01010111",
    3556 => "01010111",
    3557 => "01010111",
    3558 => "01010111",
    3559 => "01010111",
    3560 => "01010111",
    3561 => "01010111",
    3562 => "01010111",
    3563 => "01010111",
    3564 => "01010111",
    3565 => "01010111",
    3566 => "01010111",
    3567 => "01010111",
    3568 => "01010111",
    3569 => "01010111",
    3570 => "01010111",
    3571 => "01010110",
    3572 => "01010110",
    3573 => "01010110",
    3574 => "01010110",
    3575 => "01010110",
    3576 => "01010110",
    3577 => "01010110",
    3578 => "01010110",
    3579 => "01010110",
    3580 => "01010110",
    3581 => "01010110",
    3582 => "01010110",
    3583 => "01010110",
    3584 => "01010110",
    3585 => "01010110",
    3586 => "01010110",
    3587 => "01010110",
    3588 => "01010110",
    3589 => "01010110",
    3590 => "01010110",
    3591 => "01010110",
    3592 => "01010110",
    3593 => "01010110",
    3594 => "01010110",
    3595 => "01010110",
    3596 => "01010110",
    3597 => "01010110",
    3598 => "01010110",
    3599 => "01010110",
    3600 => "01010110",
    3601 => "01010110",
    3602 => "01010110",
    3603 => "01010110",
    3604 => "01010110",
    3605 => "01010110",
    3606 => "01010110",
    3607 => "01010110",
    3608 => "01010110",
    3609 => "01010110",
    3610 => "01010110",
    3611 => "01010110",
    3612 => "01010110",
    3613 => "01010101",
    3614 => "01010101",
    3615 => "01010101",
    3616 => "01010101",
    3617 => "01010101",
    3618 => "01010101",
    3619 => "01010101",
    3620 => "01010101",
    3621 => "01010101",
    3622 => "01010101",
    3623 => "01010101",
    3624 => "01010101",
    3625 => "01010101",
    3626 => "01010101",
    3627 => "01010101",
    3628 => "01010101",
    3629 => "01010101",
    3630 => "01010101",
    3631 => "01010101",
    3632 => "01010101",
    3633 => "01010101",
    3634 => "01010101",
    3635 => "01010101",
    3636 => "01010101",
    3637 => "01010101",
    3638 => "01010101",
    3639 => "01010101",
    3640 => "01010101",
    3641 => "01010101",
    3642 => "01010101",
    3643 => "01010101",
    3644 => "01010101",
    3645 => "01010101",
    3646 => "01010101",
    3647 => "01010101",
    3648 => "01010101",
    3649 => "01010101",
    3650 => "01010101",
    3651 => "01010101",
    3652 => "01010101",
    3653 => "01010101",
    3654 => "01010101",
    3655 => "01010101",
    3656 => "01010100",
    3657 => "01010100",
    3658 => "01010100",
    3659 => "01010100",
    3660 => "01010100",
    3661 => "01010100",
    3662 => "01010100",
    3663 => "01010100",
    3664 => "01010100",
    3665 => "01010100",
    3666 => "01010100",
    3667 => "01010100",
    3668 => "01010100",
    3669 => "01010100",
    3670 => "01010100",
    3671 => "01010100",
    3672 => "01010100",
    3673 => "01010100",
    3674 => "01010100",
    3675 => "01010100",
    3676 => "01010100",
    3677 => "01010100",
    3678 => "01010100",
    3679 => "01010100",
    3680 => "01010100",
    3681 => "01010100",
    3682 => "01010100",
    3683 => "01010100",
    3684 => "01010100",
    3685 => "01010100",
    3686 => "01010100",
    3687 => "01010100",
    3688 => "01010100",
    3689 => "01010100",
    3690 => "01010100",
    3691 => "01010100",
    3692 => "01010100",
    3693 => "01010100",
    3694 => "01010100",
    3695 => "01010100",
    3696 => "01010100",
    3697 => "01010100",
    3698 => "01010011",
    3699 => "01010011",
    3700 => "01010011",
    3701 => "01010011",
    3702 => "01010011",
    3703 => "01010011",
    3704 => "01010011",
    3705 => "01010011",
    3706 => "01010011",
    3707 => "01010011",
    3708 => "01010011",
    3709 => "01010011",
    3710 => "01010011",
    3711 => "01010011",
    3712 => "01010011",
    3713 => "01010011",
    3714 => "01010011",
    3715 => "01010011",
    3716 => "01010011",
    3717 => "01010011",
    3718 => "01010011",
    3719 => "01010011",
    3720 => "01010011",
    3721 => "01010011",
    3722 => "01010011",
    3723 => "01010011",
    3724 => "01010011",
    3725 => "01010011",
    3726 => "01010011",
    3727 => "01010011",
    3728 => "01010011",
    3729 => "01010011",
    3730 => "01010011",
    3731 => "01010011",
    3732 => "01010011",
    3733 => "01010011",
    3734 => "01010011",
    3735 => "01010011",
    3736 => "01010011",
    3737 => "01010011",
    3738 => "01010011",
    3739 => "01010011",
    3740 => "01010011",
    3741 => "01010011",
    3742 => "01010010",
    3743 => "01010010",
    3744 => "01010010",
    3745 => "01010010",
    3746 => "01010010",
    3747 => "01010010",
    3748 => "01010010",
    3749 => "01010010",
    3750 => "01010010",
    3751 => "01010010",
    3752 => "01010010",
    3753 => "01010010",
    3754 => "01010010",
    3755 => "01010010",
    3756 => "01010010",
    3757 => "01010010",
    3758 => "01010010",
    3759 => "01010010",
    3760 => "01010010",
    3761 => "01010010",
    3762 => "01010010",
    3763 => "01010010",
    3764 => "01010010",
    3765 => "01010010",
    3766 => "01010010",
    3767 => "01010010",
    3768 => "01010010",
    3769 => "01010010",
    3770 => "01010010",
    3771 => "01010010",
    3772 => "01010010",
    3773 => "01010010",
    3774 => "01010010",
    3775 => "01010010",
    3776 => "01010010",
    3777 => "01010010",
    3778 => "01010010",
    3779 => "01010010",
    3780 => "01010010",
    3781 => "01010010",
    3782 => "01010010",
    3783 => "01010010",
    3784 => "01010010",
    3785 => "01010001",
    3786 => "01010001",
    3787 => "01010001",
    3788 => "01010001",
    3789 => "01010001",
    3790 => "01010001",
    3791 => "01010001",
    3792 => "01010001",
    3793 => "01010001",
    3794 => "01010001",
    3795 => "01010001",
    3796 => "01010001",
    3797 => "01010001",
    3798 => "01010001",
    3799 => "01010001",
    3800 => "01010001",
    3801 => "01010001",
    3802 => "01010001",
    3803 => "01010001",
    3804 => "01010001",
    3805 => "01010001",
    3806 => "01010001",
    3807 => "01010001",
    3808 => "01010001",
    3809 => "01010001",
    3810 => "01010001",
    3811 => "01010001",
    3812 => "01010001",
    3813 => "01010001",
    3814 => "01010001",
    3815 => "01010001",
    3816 => "01010001",
    3817 => "01010001",
    3818 => "01010001",
    3819 => "01010001",
    3820 => "01010001",
    3821 => "01010001",
    3822 => "01010001",
    3823 => "01010001",
    3824 => "01010001",
    3825 => "01010001",
    3826 => "01010001",
    3827 => "01010001",
    3828 => "01010001",
    3829 => "01010000",
    3830 => "01010000",
    3831 => "01010000",
    3832 => "01010000",
    3833 => "01010000",
    3834 => "01010000",
    3835 => "01010000",
    3836 => "01010000",
    3837 => "01010000",
    3838 => "01010000",
    3839 => "01010000",
    3840 => "01010000",
    3841 => "01010000",
    3842 => "01010000",
    3843 => "01010000",
    3844 => "01010000",
    3845 => "01010000",
    3846 => "01010000",
    3847 => "01010000",
    3848 => "01010000",
    3849 => "01010000",
    3850 => "01010000",
    3851 => "01010000",
    3852 => "01010000",
    3853 => "01010000",
    3854 => "01010000",
    3855 => "01010000",
    3856 => "01010000",
    3857 => "01010000",
    3858 => "01010000",
    3859 => "01010000",
    3860 => "01010000",
    3861 => "01010000",
    3862 => "01010000",
    3863 => "01010000",
    3864 => "01010000",
    3865 => "01010000",
    3866 => "01010000",
    3867 => "01010000",
    3868 => "01010000",
    3869 => "01010000",
    3870 => "01010000",
    3871 => "01010000",
    3872 => "01001111",
    3873 => "01001111",
    3874 => "01001111",
    3875 => "01001111",
    3876 => "01001111",
    3877 => "01001111",
    3878 => "01001111",
    3879 => "01001111",
    3880 => "01001111",
    3881 => "01001111",
    3882 => "01001111",
    3883 => "01001111",
    3884 => "01001111",
    3885 => "01001111",
    3886 => "01001111",
    3887 => "01001111",
    3888 => "01001111",
    3889 => "01001111",
    3890 => "01001111",
    3891 => "01001111",
    3892 => "01001111",
    3893 => "01001111",
    3894 => "01001111",
    3895 => "01001111",
    3896 => "01001111",
    3897 => "01001111",
    3898 => "01001111",
    3899 => "01001111",
    3900 => "01001111",
    3901 => "01001111",
    3902 => "01001111",
    3903 => "01001111",
    3904 => "01001111",
    3905 => "01001111",
    3906 => "01001111",
    3907 => "01001111",
    3908 => "01001111",
    3909 => "01001111",
    3910 => "01001111",
    3911 => "01001111",
    3912 => "01001111",
    3913 => "01001111",
    3914 => "01001111",
    3915 => "01001111",
    3916 => "01001111",
    3917 => "01001110",
    3918 => "01001110",
    3919 => "01001110",
    3920 => "01001110",
    3921 => "01001110",
    3922 => "01001110",
    3923 => "01001110",
    3924 => "01001110",
    3925 => "01001110",
    3926 => "01001110",
    3927 => "01001110",
    3928 => "01001110",
    3929 => "01001110",
    3930 => "01001110",
    3931 => "01001110",
    3932 => "01001110",
    3933 => "01001110",
    3934 => "01001110",
    3935 => "01001110",
    3936 => "01001110",
    3937 => "01001110",
    3938 => "01001110",
    3939 => "01001110",
    3940 => "01001110",
    3941 => "01001110",
    3942 => "01001110",
    3943 => "01001110",
    3944 => "01001110",
    3945 => "01001110",
    3946 => "01001110",
    3947 => "01001110",
    3948 => "01001110",
    3949 => "01001110",
    3950 => "01001110",
    3951 => "01001110",
    3952 => "01001110",
    3953 => "01001110",
    3954 => "01001110",
    3955 => "01001110",
    3956 => "01001110",
    3957 => "01001110",
    3958 => "01001110",
    3959 => "01001110",
    3960 => "01001110",
    3961 => "01001101",
    3962 => "01001101",
    3963 => "01001101",
    3964 => "01001101",
    3965 => "01001101",
    3966 => "01001101",
    3967 => "01001101",
    3968 => "01001101",
    3969 => "01001101",
    3970 => "01001101",
    3971 => "01001101",
    3972 => "01001101",
    3973 => "01001101",
    3974 => "01001101",
    3975 => "01001101",
    3976 => "01001101",
    3977 => "01001101",
    3978 => "01001101",
    3979 => "01001101",
    3980 => "01001101",
    3981 => "01001101",
    3982 => "01001101",
    3983 => "01001101",
    3984 => "01001101",
    3985 => "01001101",
    3986 => "01001101",
    3987 => "01001101",
    3988 => "01001101",
    3989 => "01001101",
    3990 => "01001101",
    3991 => "01001101",
    3992 => "01001101",
    3993 => "01001101",
    3994 => "01001101",
    3995 => "01001101",
    3996 => "01001101",
    3997 => "01001101",
    3998 => "01001101",
    3999 => "01001101",
    4000 => "01001101",
    4001 => "01001101",
    4002 => "01001101",
    4003 => "01001101",
    4004 => "01001101",
    4005 => "01001101",
    4006 => "01001100",
    4007 => "01001100",
    4008 => "01001100",
    4009 => "01001100",
    4010 => "01001100",
    4011 => "01001100",
    4012 => "01001100",
    4013 => "01001100",
    4014 => "01001100",
    4015 => "01001100",
    4016 => "01001100",
    4017 => "01001100",
    4018 => "01001100",
    4019 => "01001100",
    4020 => "01001100",
    4021 => "01001100",
    4022 => "01001100",
    4023 => "01001100",
    4024 => "01001100",
    4025 => "01001100",
    4026 => "01001100",
    4027 => "01001100",
    4028 => "01001100",
    4029 => "01001100",
    4030 => "01001100",
    4031 => "01001100",
    4032 => "01001100",
    4033 => "01001100",
    4034 => "01001100",
    4035 => "01001100",
    4036 => "01001100",
    4037 => "01001100",
    4038 => "01001100",
    4039 => "01001100",
    4040 => "01001100",
    4041 => "01001100",
    4042 => "01001100",
    4043 => "01001100",
    4044 => "01001100",
    4045 => "01001100",
    4046 => "01001100",
    4047 => "01001100",
    4048 => "01001100",
    4049 => "01001100",
    4050 => "01001011",
    4051 => "01001011",
    4052 => "01001011",
    4053 => "01001011",
    4054 => "01001011",
    4055 => "01001011",
    4056 => "01001011",
    4057 => "01001011",
    4058 => "01001011",
    4059 => "01001011",
    4060 => "01001011",
    4061 => "01001011",
    4062 => "01001011",
    4063 => "01001011",
    4064 => "01001011",
    4065 => "01001011",
    4066 => "01001011",
    4067 => "01001011",
    4068 => "01001011",
    4069 => "01001011",
    4070 => "01001011",
    4071 => "01001011",
    4072 => "01001011",
    4073 => "01001011",
    4074 => "01001011",
    4075 => "01001011",
    4076 => "01001011",
    4077 => "01001011",
    4078 => "01001011",
    4079 => "01001011",
    4080 => "01001011",
    4081 => "01001011",
    4082 => "01001011",
    4083 => "01001011",
    4084 => "01001011",
    4085 => "01001011",
    4086 => "01001011",
    4087 => "01001011",
    4088 => "01001011",
    4089 => "01001011",
    4090 => "01001011",
    4091 => "01001011",
    4092 => "01001011",
    4093 => "01001011",
    4094 => "01001011",
    4095 => "01001011");
  signal q_unbuf : std_logic_vector(7 downto 0);
begin
   process (address)
   begin
     case address is
      when "000000000000" => q_unbuf <= my_rom(0);
      when "000000000001" => q_unbuf <= my_rom(1);
      when "000000000010" => q_unbuf <= my_rom(2);
      when "000000000011" => q_unbuf <= my_rom(3);
      when "000000000100" => q_unbuf <= my_rom(4);
      when "000000000101" => q_unbuf <= my_rom(5);
      when "000000000110" => q_unbuf <= my_rom(6);
      when "000000000111" => q_unbuf <= my_rom(7);
      when "000000001000" => q_unbuf <= my_rom(8);
      when "000000001001" => q_unbuf <= my_rom(9);
      when "000000001010" => q_unbuf <= my_rom(10);
      when "000000001011" => q_unbuf <= my_rom(11);
      when "000000001100" => q_unbuf <= my_rom(12);
      when "000000001101" => q_unbuf <= my_rom(13);
      when "000000001110" => q_unbuf <= my_rom(14);
      when "000000001111" => q_unbuf <= my_rom(15);
      when "000000010000" => q_unbuf <= my_rom(16);
      when "000000010001" => q_unbuf <= my_rom(17);
      when "000000010010" => q_unbuf <= my_rom(18);
      when "000000010011" => q_unbuf <= my_rom(19);
      when "000000010100" => q_unbuf <= my_rom(20);
      when "000000010101" => q_unbuf <= my_rom(21);
      when "000000010110" => q_unbuf <= my_rom(22);
      when "000000010111" => q_unbuf <= my_rom(23);
      when "000000011000" => q_unbuf <= my_rom(24);
      when "000000011001" => q_unbuf <= my_rom(25);
      when "000000011010" => q_unbuf <= my_rom(26);
      when "000000011011" => q_unbuf <= my_rom(27);
      when "000000011100" => q_unbuf <= my_rom(28);
      when "000000011101" => q_unbuf <= my_rom(29);
      when "000000011110" => q_unbuf <= my_rom(30);
      when "000000011111" => q_unbuf <= my_rom(31);
      when "000000100000" => q_unbuf <= my_rom(32);
      when "000000100001" => q_unbuf <= my_rom(33);
      when "000000100010" => q_unbuf <= my_rom(34);
      when "000000100011" => q_unbuf <= my_rom(35);
      when "000000100100" => q_unbuf <= my_rom(36);
      when "000000100101" => q_unbuf <= my_rom(37);
      when "000000100110" => q_unbuf <= my_rom(38);
      when "000000100111" => q_unbuf <= my_rom(39);
      when "000000101000" => q_unbuf <= my_rom(40);
      when "000000101001" => q_unbuf <= my_rom(41);
      when "000000101010" => q_unbuf <= my_rom(42);
      when "000000101011" => q_unbuf <= my_rom(43);
      when "000000101100" => q_unbuf <= my_rom(44);
      when "000000101101" => q_unbuf <= my_rom(45);
      when "000000101110" => q_unbuf <= my_rom(46);
      when "000000101111" => q_unbuf <= my_rom(47);
      when "000000110000" => q_unbuf <= my_rom(48);
      when "000000110001" => q_unbuf <= my_rom(49);
      when "000000110010" => q_unbuf <= my_rom(50);
      when "000000110011" => q_unbuf <= my_rom(51);
      when "000000110100" => q_unbuf <= my_rom(52);
      when "000000110101" => q_unbuf <= my_rom(53);
      when "000000110110" => q_unbuf <= my_rom(54);
      when "000000110111" => q_unbuf <= my_rom(55);
      when "000000111000" => q_unbuf <= my_rom(56);
      when "000000111001" => q_unbuf <= my_rom(57);
      when "000000111010" => q_unbuf <= my_rom(58);
      when "000000111011" => q_unbuf <= my_rom(59);
      when "000000111100" => q_unbuf <= my_rom(60);
      when "000000111101" => q_unbuf <= my_rom(61);
      when "000000111110" => q_unbuf <= my_rom(62);
      when "000000111111" => q_unbuf <= my_rom(63);
      when "000001000000" => q_unbuf <= my_rom(64);
      when "000001000001" => q_unbuf <= my_rom(65);
      when "000001000010" => q_unbuf <= my_rom(66);
      when "000001000011" => q_unbuf <= my_rom(67);
      when "000001000100" => q_unbuf <= my_rom(68);
      when "000001000101" => q_unbuf <= my_rom(69);
      when "000001000110" => q_unbuf <= my_rom(70);
      when "000001000111" => q_unbuf <= my_rom(71);
      when "000001001000" => q_unbuf <= my_rom(72);
      when "000001001001" => q_unbuf <= my_rom(73);
      when "000001001010" => q_unbuf <= my_rom(74);
      when "000001001011" => q_unbuf <= my_rom(75);
      when "000001001100" => q_unbuf <= my_rom(76);
      when "000001001101" => q_unbuf <= my_rom(77);
      when "000001001110" => q_unbuf <= my_rom(78);
      when "000001001111" => q_unbuf <= my_rom(79);
      when "000001010000" => q_unbuf <= my_rom(80);
      when "000001010001" => q_unbuf <= my_rom(81);
      when "000001010010" => q_unbuf <= my_rom(82);
      when "000001010011" => q_unbuf <= my_rom(83);
      when "000001010100" => q_unbuf <= my_rom(84);
      when "000001010101" => q_unbuf <= my_rom(85);
      when "000001010110" => q_unbuf <= my_rom(86);
      when "000001010111" => q_unbuf <= my_rom(87);
      when "000001011000" => q_unbuf <= my_rom(88);
      when "000001011001" => q_unbuf <= my_rom(89);
      when "000001011010" => q_unbuf <= my_rom(90);
      when "000001011011" => q_unbuf <= my_rom(91);
      when "000001011100" => q_unbuf <= my_rom(92);
      when "000001011101" => q_unbuf <= my_rom(93);
      when "000001011110" => q_unbuf <= my_rom(94);
      when "000001011111" => q_unbuf <= my_rom(95);
      when "000001100000" => q_unbuf <= my_rom(96);
      when "000001100001" => q_unbuf <= my_rom(97);
      when "000001100010" => q_unbuf <= my_rom(98);
      when "000001100011" => q_unbuf <= my_rom(99);
      when "000001100100" => q_unbuf <= my_rom(100);
      when "000001100101" => q_unbuf <= my_rom(101);
      when "000001100110" => q_unbuf <= my_rom(102);
      when "000001100111" => q_unbuf <= my_rom(103);
      when "000001101000" => q_unbuf <= my_rom(104);
      when "000001101001" => q_unbuf <= my_rom(105);
      when "000001101010" => q_unbuf <= my_rom(106);
      when "000001101011" => q_unbuf <= my_rom(107);
      when "000001101100" => q_unbuf <= my_rom(108);
      when "000001101101" => q_unbuf <= my_rom(109);
      when "000001101110" => q_unbuf <= my_rom(110);
      when "000001101111" => q_unbuf <= my_rom(111);
      when "000001110000" => q_unbuf <= my_rom(112);
      when "000001110001" => q_unbuf <= my_rom(113);
      when "000001110010" => q_unbuf <= my_rom(114);
      when "000001110011" => q_unbuf <= my_rom(115);
      when "000001110100" => q_unbuf <= my_rom(116);
      when "000001110101" => q_unbuf <= my_rom(117);
      when "000001110110" => q_unbuf <= my_rom(118);
      when "000001110111" => q_unbuf <= my_rom(119);
      when "000001111000" => q_unbuf <= my_rom(120);
      when "000001111001" => q_unbuf <= my_rom(121);
      when "000001111010" => q_unbuf <= my_rom(122);
      when "000001111011" => q_unbuf <= my_rom(123);
      when "000001111100" => q_unbuf <= my_rom(124);
      when "000001111101" => q_unbuf <= my_rom(125);
      when "000001111110" => q_unbuf <= my_rom(126);
      when "000001111111" => q_unbuf <= my_rom(127);
      when "000010000000" => q_unbuf <= my_rom(128);
      when "000010000001" => q_unbuf <= my_rom(129);
      when "000010000010" => q_unbuf <= my_rom(130);
      when "000010000011" => q_unbuf <= my_rom(131);
      when "000010000100" => q_unbuf <= my_rom(132);
      when "000010000101" => q_unbuf <= my_rom(133);
      when "000010000110" => q_unbuf <= my_rom(134);
      when "000010000111" => q_unbuf <= my_rom(135);
      when "000010001000" => q_unbuf <= my_rom(136);
      when "000010001001" => q_unbuf <= my_rom(137);
      when "000010001010" => q_unbuf <= my_rom(138);
      when "000010001011" => q_unbuf <= my_rom(139);
      when "000010001100" => q_unbuf <= my_rom(140);
      when "000010001101" => q_unbuf <= my_rom(141);
      when "000010001110" => q_unbuf <= my_rom(142);
      when "000010001111" => q_unbuf <= my_rom(143);
      when "000010010000" => q_unbuf <= my_rom(144);
      when "000010010001" => q_unbuf <= my_rom(145);
      when "000010010010" => q_unbuf <= my_rom(146);
      when "000010010011" => q_unbuf <= my_rom(147);
      when "000010010100" => q_unbuf <= my_rom(148);
      when "000010010101" => q_unbuf <= my_rom(149);
      when "000010010110" => q_unbuf <= my_rom(150);
      when "000010010111" => q_unbuf <= my_rom(151);
      when "000010011000" => q_unbuf <= my_rom(152);
      when "000010011001" => q_unbuf <= my_rom(153);
      when "000010011010" => q_unbuf <= my_rom(154);
      when "000010011011" => q_unbuf <= my_rom(155);
      when "000010011100" => q_unbuf <= my_rom(156);
      when "000010011101" => q_unbuf <= my_rom(157);
      when "000010011110" => q_unbuf <= my_rom(158);
      when "000010011111" => q_unbuf <= my_rom(159);
      when "000010100000" => q_unbuf <= my_rom(160);
      when "000010100001" => q_unbuf <= my_rom(161);
      when "000010100010" => q_unbuf <= my_rom(162);
      when "000010100011" => q_unbuf <= my_rom(163);
      when "000010100100" => q_unbuf <= my_rom(164);
      when "000010100101" => q_unbuf <= my_rom(165);
      when "000010100110" => q_unbuf <= my_rom(166);
      when "000010100111" => q_unbuf <= my_rom(167);
      when "000010101000" => q_unbuf <= my_rom(168);
      when "000010101001" => q_unbuf <= my_rom(169);
      when "000010101010" => q_unbuf <= my_rom(170);
      when "000010101011" => q_unbuf <= my_rom(171);
      when "000010101100" => q_unbuf <= my_rom(172);
      when "000010101101" => q_unbuf <= my_rom(173);
      when "000010101110" => q_unbuf <= my_rom(174);
      when "000010101111" => q_unbuf <= my_rom(175);
      when "000010110000" => q_unbuf <= my_rom(176);
      when "000010110001" => q_unbuf <= my_rom(177);
      when "000010110010" => q_unbuf <= my_rom(178);
      when "000010110011" => q_unbuf <= my_rom(179);
      when "000010110100" => q_unbuf <= my_rom(180);
      when "000010110101" => q_unbuf <= my_rom(181);
      when "000010110110" => q_unbuf <= my_rom(182);
      when "000010110111" => q_unbuf <= my_rom(183);
      when "000010111000" => q_unbuf <= my_rom(184);
      when "000010111001" => q_unbuf <= my_rom(185);
      when "000010111010" => q_unbuf <= my_rom(186);
      when "000010111011" => q_unbuf <= my_rom(187);
      when "000010111100" => q_unbuf <= my_rom(188);
      when "000010111101" => q_unbuf <= my_rom(189);
      when "000010111110" => q_unbuf <= my_rom(190);
      when "000010111111" => q_unbuf <= my_rom(191);
      when "000011000000" => q_unbuf <= my_rom(192);
      when "000011000001" => q_unbuf <= my_rom(193);
      when "000011000010" => q_unbuf <= my_rom(194);
      when "000011000011" => q_unbuf <= my_rom(195);
      when "000011000100" => q_unbuf <= my_rom(196);
      when "000011000101" => q_unbuf <= my_rom(197);
      when "000011000110" => q_unbuf <= my_rom(198);
      when "000011000111" => q_unbuf <= my_rom(199);
      when "000011001000" => q_unbuf <= my_rom(200);
      when "000011001001" => q_unbuf <= my_rom(201);
      when "000011001010" => q_unbuf <= my_rom(202);
      when "000011001011" => q_unbuf <= my_rom(203);
      when "000011001100" => q_unbuf <= my_rom(204);
      when "000011001101" => q_unbuf <= my_rom(205);
      when "000011001110" => q_unbuf <= my_rom(206);
      when "000011001111" => q_unbuf <= my_rom(207);
      when "000011010000" => q_unbuf <= my_rom(208);
      when "000011010001" => q_unbuf <= my_rom(209);
      when "000011010010" => q_unbuf <= my_rom(210);
      when "000011010011" => q_unbuf <= my_rom(211);
      when "000011010100" => q_unbuf <= my_rom(212);
      when "000011010101" => q_unbuf <= my_rom(213);
      when "000011010110" => q_unbuf <= my_rom(214);
      when "000011010111" => q_unbuf <= my_rom(215);
      when "000011011000" => q_unbuf <= my_rom(216);
      when "000011011001" => q_unbuf <= my_rom(217);
      when "000011011010" => q_unbuf <= my_rom(218);
      when "000011011011" => q_unbuf <= my_rom(219);
      when "000011011100" => q_unbuf <= my_rom(220);
      when "000011011101" => q_unbuf <= my_rom(221);
      when "000011011110" => q_unbuf <= my_rom(222);
      when "000011011111" => q_unbuf <= my_rom(223);
      when "000011100000" => q_unbuf <= my_rom(224);
      when "000011100001" => q_unbuf <= my_rom(225);
      when "000011100010" => q_unbuf <= my_rom(226);
      when "000011100011" => q_unbuf <= my_rom(227);
      when "000011100100" => q_unbuf <= my_rom(228);
      when "000011100101" => q_unbuf <= my_rom(229);
      when "000011100110" => q_unbuf <= my_rom(230);
      when "000011100111" => q_unbuf <= my_rom(231);
      when "000011101000" => q_unbuf <= my_rom(232);
      when "000011101001" => q_unbuf <= my_rom(233);
      when "000011101010" => q_unbuf <= my_rom(234);
      when "000011101011" => q_unbuf <= my_rom(235);
      when "000011101100" => q_unbuf <= my_rom(236);
      when "000011101101" => q_unbuf <= my_rom(237);
      when "000011101110" => q_unbuf <= my_rom(238);
      when "000011101111" => q_unbuf <= my_rom(239);
      when "000011110000" => q_unbuf <= my_rom(240);
      when "000011110001" => q_unbuf <= my_rom(241);
      when "000011110010" => q_unbuf <= my_rom(242);
      when "000011110011" => q_unbuf <= my_rom(243);
      when "000011110100" => q_unbuf <= my_rom(244);
      when "000011110101" => q_unbuf <= my_rom(245);
      when "000011110110" => q_unbuf <= my_rom(246);
      when "000011110111" => q_unbuf <= my_rom(247);
      when "000011111000" => q_unbuf <= my_rom(248);
      when "000011111001" => q_unbuf <= my_rom(249);
      when "000011111010" => q_unbuf <= my_rom(250);
      when "000011111011" => q_unbuf <= my_rom(251);
      when "000011111100" => q_unbuf <= my_rom(252);
      when "000011111101" => q_unbuf <= my_rom(253);
      when "000011111110" => q_unbuf <= my_rom(254);
      when "000011111111" => q_unbuf <= my_rom(255);
      when "000100000000" => q_unbuf <= my_rom(256);
      when "000100000001" => q_unbuf <= my_rom(257);
      when "000100000010" => q_unbuf <= my_rom(258);
      when "000100000011" => q_unbuf <= my_rom(259);
      when "000100000100" => q_unbuf <= my_rom(260);
      when "000100000101" => q_unbuf <= my_rom(261);
      when "000100000110" => q_unbuf <= my_rom(262);
      when "000100000111" => q_unbuf <= my_rom(263);
      when "000100001000" => q_unbuf <= my_rom(264);
      when "000100001001" => q_unbuf <= my_rom(265);
      when "000100001010" => q_unbuf <= my_rom(266);
      when "000100001011" => q_unbuf <= my_rom(267);
      when "000100001100" => q_unbuf <= my_rom(268);
      when "000100001101" => q_unbuf <= my_rom(269);
      when "000100001110" => q_unbuf <= my_rom(270);
      when "000100001111" => q_unbuf <= my_rom(271);
      when "000100010000" => q_unbuf <= my_rom(272);
      when "000100010001" => q_unbuf <= my_rom(273);
      when "000100010010" => q_unbuf <= my_rom(274);
      when "000100010011" => q_unbuf <= my_rom(275);
      when "000100010100" => q_unbuf <= my_rom(276);
      when "000100010101" => q_unbuf <= my_rom(277);
      when "000100010110" => q_unbuf <= my_rom(278);
      when "000100010111" => q_unbuf <= my_rom(279);
      when "000100011000" => q_unbuf <= my_rom(280);
      when "000100011001" => q_unbuf <= my_rom(281);
      when "000100011010" => q_unbuf <= my_rom(282);
      when "000100011011" => q_unbuf <= my_rom(283);
      when "000100011100" => q_unbuf <= my_rom(284);
      when "000100011101" => q_unbuf <= my_rom(285);
      when "000100011110" => q_unbuf <= my_rom(286);
      when "000100011111" => q_unbuf <= my_rom(287);
      when "000100100000" => q_unbuf <= my_rom(288);
      when "000100100001" => q_unbuf <= my_rom(289);
      when "000100100010" => q_unbuf <= my_rom(290);
      when "000100100011" => q_unbuf <= my_rom(291);
      when "000100100100" => q_unbuf <= my_rom(292);
      when "000100100101" => q_unbuf <= my_rom(293);
      when "000100100110" => q_unbuf <= my_rom(294);
      when "000100100111" => q_unbuf <= my_rom(295);
      when "000100101000" => q_unbuf <= my_rom(296);
      when "000100101001" => q_unbuf <= my_rom(297);
      when "000100101010" => q_unbuf <= my_rom(298);
      when "000100101011" => q_unbuf <= my_rom(299);
      when "000100101100" => q_unbuf <= my_rom(300);
      when "000100101101" => q_unbuf <= my_rom(301);
      when "000100101110" => q_unbuf <= my_rom(302);
      when "000100101111" => q_unbuf <= my_rom(303);
      when "000100110000" => q_unbuf <= my_rom(304);
      when "000100110001" => q_unbuf <= my_rom(305);
      when "000100110010" => q_unbuf <= my_rom(306);
      when "000100110011" => q_unbuf <= my_rom(307);
      when "000100110100" => q_unbuf <= my_rom(308);
      when "000100110101" => q_unbuf <= my_rom(309);
      when "000100110110" => q_unbuf <= my_rom(310);
      when "000100110111" => q_unbuf <= my_rom(311);
      when "000100111000" => q_unbuf <= my_rom(312);
      when "000100111001" => q_unbuf <= my_rom(313);
      when "000100111010" => q_unbuf <= my_rom(314);
      when "000100111011" => q_unbuf <= my_rom(315);
      when "000100111100" => q_unbuf <= my_rom(316);
      when "000100111101" => q_unbuf <= my_rom(317);
      when "000100111110" => q_unbuf <= my_rom(318);
      when "000100111111" => q_unbuf <= my_rom(319);
      when "000101000000" => q_unbuf <= my_rom(320);
      when "000101000001" => q_unbuf <= my_rom(321);
      when "000101000010" => q_unbuf <= my_rom(322);
      when "000101000011" => q_unbuf <= my_rom(323);
      when "000101000100" => q_unbuf <= my_rom(324);
      when "000101000101" => q_unbuf <= my_rom(325);
      when "000101000110" => q_unbuf <= my_rom(326);
      when "000101000111" => q_unbuf <= my_rom(327);
      when "000101001000" => q_unbuf <= my_rom(328);
      when "000101001001" => q_unbuf <= my_rom(329);
      when "000101001010" => q_unbuf <= my_rom(330);
      when "000101001011" => q_unbuf <= my_rom(331);
      when "000101001100" => q_unbuf <= my_rom(332);
      when "000101001101" => q_unbuf <= my_rom(333);
      when "000101001110" => q_unbuf <= my_rom(334);
      when "000101001111" => q_unbuf <= my_rom(335);
      when "000101010000" => q_unbuf <= my_rom(336);
      when "000101010001" => q_unbuf <= my_rom(337);
      when "000101010010" => q_unbuf <= my_rom(338);
      when "000101010011" => q_unbuf <= my_rom(339);
      when "000101010100" => q_unbuf <= my_rom(340);
      when "000101010101" => q_unbuf <= my_rom(341);
      when "000101010110" => q_unbuf <= my_rom(342);
      when "000101010111" => q_unbuf <= my_rom(343);
      when "000101011000" => q_unbuf <= my_rom(344);
      when "000101011001" => q_unbuf <= my_rom(345);
      when "000101011010" => q_unbuf <= my_rom(346);
      when "000101011011" => q_unbuf <= my_rom(347);
      when "000101011100" => q_unbuf <= my_rom(348);
      when "000101011101" => q_unbuf <= my_rom(349);
      when "000101011110" => q_unbuf <= my_rom(350);
      when "000101011111" => q_unbuf <= my_rom(351);
      when "000101100000" => q_unbuf <= my_rom(352);
      when "000101100001" => q_unbuf <= my_rom(353);
      when "000101100010" => q_unbuf <= my_rom(354);
      when "000101100011" => q_unbuf <= my_rom(355);
      when "000101100100" => q_unbuf <= my_rom(356);
      when "000101100101" => q_unbuf <= my_rom(357);
      when "000101100110" => q_unbuf <= my_rom(358);
      when "000101100111" => q_unbuf <= my_rom(359);
      when "000101101000" => q_unbuf <= my_rom(360);
      when "000101101001" => q_unbuf <= my_rom(361);
      when "000101101010" => q_unbuf <= my_rom(362);
      when "000101101011" => q_unbuf <= my_rom(363);
      when "000101101100" => q_unbuf <= my_rom(364);
      when "000101101101" => q_unbuf <= my_rom(365);
      when "000101101110" => q_unbuf <= my_rom(366);
      when "000101101111" => q_unbuf <= my_rom(367);
      when "000101110000" => q_unbuf <= my_rom(368);
      when "000101110001" => q_unbuf <= my_rom(369);
      when "000101110010" => q_unbuf <= my_rom(370);
      when "000101110011" => q_unbuf <= my_rom(371);
      when "000101110100" => q_unbuf <= my_rom(372);
      when "000101110101" => q_unbuf <= my_rom(373);
      when "000101110110" => q_unbuf <= my_rom(374);
      when "000101110111" => q_unbuf <= my_rom(375);
      when "000101111000" => q_unbuf <= my_rom(376);
      when "000101111001" => q_unbuf <= my_rom(377);
      when "000101111010" => q_unbuf <= my_rom(378);
      when "000101111011" => q_unbuf <= my_rom(379);
      when "000101111100" => q_unbuf <= my_rom(380);
      when "000101111101" => q_unbuf <= my_rom(381);
      when "000101111110" => q_unbuf <= my_rom(382);
      when "000101111111" => q_unbuf <= my_rom(383);
      when "000110000000" => q_unbuf <= my_rom(384);
      when "000110000001" => q_unbuf <= my_rom(385);
      when "000110000010" => q_unbuf <= my_rom(386);
      when "000110000011" => q_unbuf <= my_rom(387);
      when "000110000100" => q_unbuf <= my_rom(388);
      when "000110000101" => q_unbuf <= my_rom(389);
      when "000110000110" => q_unbuf <= my_rom(390);
      when "000110000111" => q_unbuf <= my_rom(391);
      when "000110001000" => q_unbuf <= my_rom(392);
      when "000110001001" => q_unbuf <= my_rom(393);
      when "000110001010" => q_unbuf <= my_rom(394);
      when "000110001011" => q_unbuf <= my_rom(395);
      when "000110001100" => q_unbuf <= my_rom(396);
      when "000110001101" => q_unbuf <= my_rom(397);
      when "000110001110" => q_unbuf <= my_rom(398);
      when "000110001111" => q_unbuf <= my_rom(399);
      when "000110010000" => q_unbuf <= my_rom(400);
      when "000110010001" => q_unbuf <= my_rom(401);
      when "000110010010" => q_unbuf <= my_rom(402);
      when "000110010011" => q_unbuf <= my_rom(403);
      when "000110010100" => q_unbuf <= my_rom(404);
      when "000110010101" => q_unbuf <= my_rom(405);
      when "000110010110" => q_unbuf <= my_rom(406);
      when "000110010111" => q_unbuf <= my_rom(407);
      when "000110011000" => q_unbuf <= my_rom(408);
      when "000110011001" => q_unbuf <= my_rom(409);
      when "000110011010" => q_unbuf <= my_rom(410);
      when "000110011011" => q_unbuf <= my_rom(411);
      when "000110011100" => q_unbuf <= my_rom(412);
      when "000110011101" => q_unbuf <= my_rom(413);
      when "000110011110" => q_unbuf <= my_rom(414);
      when "000110011111" => q_unbuf <= my_rom(415);
      when "000110100000" => q_unbuf <= my_rom(416);
      when "000110100001" => q_unbuf <= my_rom(417);
      when "000110100010" => q_unbuf <= my_rom(418);
      when "000110100011" => q_unbuf <= my_rom(419);
      when "000110100100" => q_unbuf <= my_rom(420);
      when "000110100101" => q_unbuf <= my_rom(421);
      when "000110100110" => q_unbuf <= my_rom(422);
      when "000110100111" => q_unbuf <= my_rom(423);
      when "000110101000" => q_unbuf <= my_rom(424);
      when "000110101001" => q_unbuf <= my_rom(425);
      when "000110101010" => q_unbuf <= my_rom(426);
      when "000110101011" => q_unbuf <= my_rom(427);
      when "000110101100" => q_unbuf <= my_rom(428);
      when "000110101101" => q_unbuf <= my_rom(429);
      when "000110101110" => q_unbuf <= my_rom(430);
      when "000110101111" => q_unbuf <= my_rom(431);
      when "000110110000" => q_unbuf <= my_rom(432);
      when "000110110001" => q_unbuf <= my_rom(433);
      when "000110110010" => q_unbuf <= my_rom(434);
      when "000110110011" => q_unbuf <= my_rom(435);
      when "000110110100" => q_unbuf <= my_rom(436);
      when "000110110101" => q_unbuf <= my_rom(437);
      when "000110110110" => q_unbuf <= my_rom(438);
      when "000110110111" => q_unbuf <= my_rom(439);
      when "000110111000" => q_unbuf <= my_rom(440);
      when "000110111001" => q_unbuf <= my_rom(441);
      when "000110111010" => q_unbuf <= my_rom(442);
      when "000110111011" => q_unbuf <= my_rom(443);
      when "000110111100" => q_unbuf <= my_rom(444);
      when "000110111101" => q_unbuf <= my_rom(445);
      when "000110111110" => q_unbuf <= my_rom(446);
      when "000110111111" => q_unbuf <= my_rom(447);
      when "000111000000" => q_unbuf <= my_rom(448);
      when "000111000001" => q_unbuf <= my_rom(449);
      when "000111000010" => q_unbuf <= my_rom(450);
      when "000111000011" => q_unbuf <= my_rom(451);
      when "000111000100" => q_unbuf <= my_rom(452);
      when "000111000101" => q_unbuf <= my_rom(453);
      when "000111000110" => q_unbuf <= my_rom(454);
      when "000111000111" => q_unbuf <= my_rom(455);
      when "000111001000" => q_unbuf <= my_rom(456);
      when "000111001001" => q_unbuf <= my_rom(457);
      when "000111001010" => q_unbuf <= my_rom(458);
      when "000111001011" => q_unbuf <= my_rom(459);
      when "000111001100" => q_unbuf <= my_rom(460);
      when "000111001101" => q_unbuf <= my_rom(461);
      when "000111001110" => q_unbuf <= my_rom(462);
      when "000111001111" => q_unbuf <= my_rom(463);
      when "000111010000" => q_unbuf <= my_rom(464);
      when "000111010001" => q_unbuf <= my_rom(465);
      when "000111010010" => q_unbuf <= my_rom(466);
      when "000111010011" => q_unbuf <= my_rom(467);
      when "000111010100" => q_unbuf <= my_rom(468);
      when "000111010101" => q_unbuf <= my_rom(469);
      when "000111010110" => q_unbuf <= my_rom(470);
      when "000111010111" => q_unbuf <= my_rom(471);
      when "000111011000" => q_unbuf <= my_rom(472);
      when "000111011001" => q_unbuf <= my_rom(473);
      when "000111011010" => q_unbuf <= my_rom(474);
      when "000111011011" => q_unbuf <= my_rom(475);
      when "000111011100" => q_unbuf <= my_rom(476);
      when "000111011101" => q_unbuf <= my_rom(477);
      when "000111011110" => q_unbuf <= my_rom(478);
      when "000111011111" => q_unbuf <= my_rom(479);
      when "000111100000" => q_unbuf <= my_rom(480);
      when "000111100001" => q_unbuf <= my_rom(481);
      when "000111100010" => q_unbuf <= my_rom(482);
      when "000111100011" => q_unbuf <= my_rom(483);
      when "000111100100" => q_unbuf <= my_rom(484);
      when "000111100101" => q_unbuf <= my_rom(485);
      when "000111100110" => q_unbuf <= my_rom(486);
      when "000111100111" => q_unbuf <= my_rom(487);
      when "000111101000" => q_unbuf <= my_rom(488);
      when "000111101001" => q_unbuf <= my_rom(489);
      when "000111101010" => q_unbuf <= my_rom(490);
      when "000111101011" => q_unbuf <= my_rom(491);
      when "000111101100" => q_unbuf <= my_rom(492);
      when "000111101101" => q_unbuf <= my_rom(493);
      when "000111101110" => q_unbuf <= my_rom(494);
      when "000111101111" => q_unbuf <= my_rom(495);
      when "000111110000" => q_unbuf <= my_rom(496);
      when "000111110001" => q_unbuf <= my_rom(497);
      when "000111110010" => q_unbuf <= my_rom(498);
      when "000111110011" => q_unbuf <= my_rom(499);
      when "000111110100" => q_unbuf <= my_rom(500);
      when "000111110101" => q_unbuf <= my_rom(501);
      when "000111110110" => q_unbuf <= my_rom(502);
      when "000111110111" => q_unbuf <= my_rom(503);
      when "000111111000" => q_unbuf <= my_rom(504);
      when "000111111001" => q_unbuf <= my_rom(505);
      when "000111111010" => q_unbuf <= my_rom(506);
      when "000111111011" => q_unbuf <= my_rom(507);
      when "000111111100" => q_unbuf <= my_rom(508);
      when "000111111101" => q_unbuf <= my_rom(509);
      when "000111111110" => q_unbuf <= my_rom(510);
      when "000111111111" => q_unbuf <= my_rom(511);
      when "001000000000" => q_unbuf <= my_rom(512);
      when "001000000001" => q_unbuf <= my_rom(513);
      when "001000000010" => q_unbuf <= my_rom(514);
      when "001000000011" => q_unbuf <= my_rom(515);
      when "001000000100" => q_unbuf <= my_rom(516);
      when "001000000101" => q_unbuf <= my_rom(517);
      when "001000000110" => q_unbuf <= my_rom(518);
      when "001000000111" => q_unbuf <= my_rom(519);
      when "001000001000" => q_unbuf <= my_rom(520);
      when "001000001001" => q_unbuf <= my_rom(521);
      when "001000001010" => q_unbuf <= my_rom(522);
      when "001000001011" => q_unbuf <= my_rom(523);
      when "001000001100" => q_unbuf <= my_rom(524);
      when "001000001101" => q_unbuf <= my_rom(525);
      when "001000001110" => q_unbuf <= my_rom(526);
      when "001000001111" => q_unbuf <= my_rom(527);
      when "001000010000" => q_unbuf <= my_rom(528);
      when "001000010001" => q_unbuf <= my_rom(529);
      when "001000010010" => q_unbuf <= my_rom(530);
      when "001000010011" => q_unbuf <= my_rom(531);
      when "001000010100" => q_unbuf <= my_rom(532);
      when "001000010101" => q_unbuf <= my_rom(533);
      when "001000010110" => q_unbuf <= my_rom(534);
      when "001000010111" => q_unbuf <= my_rom(535);
      when "001000011000" => q_unbuf <= my_rom(536);
      when "001000011001" => q_unbuf <= my_rom(537);
      when "001000011010" => q_unbuf <= my_rom(538);
      when "001000011011" => q_unbuf <= my_rom(539);
      when "001000011100" => q_unbuf <= my_rom(540);
      when "001000011101" => q_unbuf <= my_rom(541);
      when "001000011110" => q_unbuf <= my_rom(542);
      when "001000011111" => q_unbuf <= my_rom(543);
      when "001000100000" => q_unbuf <= my_rom(544);
      when "001000100001" => q_unbuf <= my_rom(545);
      when "001000100010" => q_unbuf <= my_rom(546);
      when "001000100011" => q_unbuf <= my_rom(547);
      when "001000100100" => q_unbuf <= my_rom(548);
      when "001000100101" => q_unbuf <= my_rom(549);
      when "001000100110" => q_unbuf <= my_rom(550);
      when "001000100111" => q_unbuf <= my_rom(551);
      when "001000101000" => q_unbuf <= my_rom(552);
      when "001000101001" => q_unbuf <= my_rom(553);
      when "001000101010" => q_unbuf <= my_rom(554);
      when "001000101011" => q_unbuf <= my_rom(555);
      when "001000101100" => q_unbuf <= my_rom(556);
      when "001000101101" => q_unbuf <= my_rom(557);
      when "001000101110" => q_unbuf <= my_rom(558);
      when "001000101111" => q_unbuf <= my_rom(559);
      when "001000110000" => q_unbuf <= my_rom(560);
      when "001000110001" => q_unbuf <= my_rom(561);
      when "001000110010" => q_unbuf <= my_rom(562);
      when "001000110011" => q_unbuf <= my_rom(563);
      when "001000110100" => q_unbuf <= my_rom(564);
      when "001000110101" => q_unbuf <= my_rom(565);
      when "001000110110" => q_unbuf <= my_rom(566);
      when "001000110111" => q_unbuf <= my_rom(567);
      when "001000111000" => q_unbuf <= my_rom(568);
      when "001000111001" => q_unbuf <= my_rom(569);
      when "001000111010" => q_unbuf <= my_rom(570);
      when "001000111011" => q_unbuf <= my_rom(571);
      when "001000111100" => q_unbuf <= my_rom(572);
      when "001000111101" => q_unbuf <= my_rom(573);
      when "001000111110" => q_unbuf <= my_rom(574);
      when "001000111111" => q_unbuf <= my_rom(575);
      when "001001000000" => q_unbuf <= my_rom(576);
      when "001001000001" => q_unbuf <= my_rom(577);
      when "001001000010" => q_unbuf <= my_rom(578);
      when "001001000011" => q_unbuf <= my_rom(579);
      when "001001000100" => q_unbuf <= my_rom(580);
      when "001001000101" => q_unbuf <= my_rom(581);
      when "001001000110" => q_unbuf <= my_rom(582);
      when "001001000111" => q_unbuf <= my_rom(583);
      when "001001001000" => q_unbuf <= my_rom(584);
      when "001001001001" => q_unbuf <= my_rom(585);
      when "001001001010" => q_unbuf <= my_rom(586);
      when "001001001011" => q_unbuf <= my_rom(587);
      when "001001001100" => q_unbuf <= my_rom(588);
      when "001001001101" => q_unbuf <= my_rom(589);
      when "001001001110" => q_unbuf <= my_rom(590);
      when "001001001111" => q_unbuf <= my_rom(591);
      when "001001010000" => q_unbuf <= my_rom(592);
      when "001001010001" => q_unbuf <= my_rom(593);
      when "001001010010" => q_unbuf <= my_rom(594);
      when "001001010011" => q_unbuf <= my_rom(595);
      when "001001010100" => q_unbuf <= my_rom(596);
      when "001001010101" => q_unbuf <= my_rom(597);
      when "001001010110" => q_unbuf <= my_rom(598);
      when "001001010111" => q_unbuf <= my_rom(599);
      when "001001011000" => q_unbuf <= my_rom(600);
      when "001001011001" => q_unbuf <= my_rom(601);
      when "001001011010" => q_unbuf <= my_rom(602);
      when "001001011011" => q_unbuf <= my_rom(603);
      when "001001011100" => q_unbuf <= my_rom(604);
      when "001001011101" => q_unbuf <= my_rom(605);
      when "001001011110" => q_unbuf <= my_rom(606);
      when "001001011111" => q_unbuf <= my_rom(607);
      when "001001100000" => q_unbuf <= my_rom(608);
      when "001001100001" => q_unbuf <= my_rom(609);
      when "001001100010" => q_unbuf <= my_rom(610);
      when "001001100011" => q_unbuf <= my_rom(611);
      when "001001100100" => q_unbuf <= my_rom(612);
      when "001001100101" => q_unbuf <= my_rom(613);
      when "001001100110" => q_unbuf <= my_rom(614);
      when "001001100111" => q_unbuf <= my_rom(615);
      when "001001101000" => q_unbuf <= my_rom(616);
      when "001001101001" => q_unbuf <= my_rom(617);
      when "001001101010" => q_unbuf <= my_rom(618);
      when "001001101011" => q_unbuf <= my_rom(619);
      when "001001101100" => q_unbuf <= my_rom(620);
      when "001001101101" => q_unbuf <= my_rom(621);
      when "001001101110" => q_unbuf <= my_rom(622);
      when "001001101111" => q_unbuf <= my_rom(623);
      when "001001110000" => q_unbuf <= my_rom(624);
      when "001001110001" => q_unbuf <= my_rom(625);
      when "001001110010" => q_unbuf <= my_rom(626);
      when "001001110011" => q_unbuf <= my_rom(627);
      when "001001110100" => q_unbuf <= my_rom(628);
      when "001001110101" => q_unbuf <= my_rom(629);
      when "001001110110" => q_unbuf <= my_rom(630);
      when "001001110111" => q_unbuf <= my_rom(631);
      when "001001111000" => q_unbuf <= my_rom(632);
      when "001001111001" => q_unbuf <= my_rom(633);
      when "001001111010" => q_unbuf <= my_rom(634);
      when "001001111011" => q_unbuf <= my_rom(635);
      when "001001111100" => q_unbuf <= my_rom(636);
      when "001001111101" => q_unbuf <= my_rom(637);
      when "001001111110" => q_unbuf <= my_rom(638);
      when "001001111111" => q_unbuf <= my_rom(639);
      when "001010000000" => q_unbuf <= my_rom(640);
      when "001010000001" => q_unbuf <= my_rom(641);
      when "001010000010" => q_unbuf <= my_rom(642);
      when "001010000011" => q_unbuf <= my_rom(643);
      when "001010000100" => q_unbuf <= my_rom(644);
      when "001010000101" => q_unbuf <= my_rom(645);
      when "001010000110" => q_unbuf <= my_rom(646);
      when "001010000111" => q_unbuf <= my_rom(647);
      when "001010001000" => q_unbuf <= my_rom(648);
      when "001010001001" => q_unbuf <= my_rom(649);
      when "001010001010" => q_unbuf <= my_rom(650);
      when "001010001011" => q_unbuf <= my_rom(651);
      when "001010001100" => q_unbuf <= my_rom(652);
      when "001010001101" => q_unbuf <= my_rom(653);
      when "001010001110" => q_unbuf <= my_rom(654);
      when "001010001111" => q_unbuf <= my_rom(655);
      when "001010010000" => q_unbuf <= my_rom(656);
      when "001010010001" => q_unbuf <= my_rom(657);
      when "001010010010" => q_unbuf <= my_rom(658);
      when "001010010011" => q_unbuf <= my_rom(659);
      when "001010010100" => q_unbuf <= my_rom(660);
      when "001010010101" => q_unbuf <= my_rom(661);
      when "001010010110" => q_unbuf <= my_rom(662);
      when "001010010111" => q_unbuf <= my_rom(663);
      when "001010011000" => q_unbuf <= my_rom(664);
      when "001010011001" => q_unbuf <= my_rom(665);
      when "001010011010" => q_unbuf <= my_rom(666);
      when "001010011011" => q_unbuf <= my_rom(667);
      when "001010011100" => q_unbuf <= my_rom(668);
      when "001010011101" => q_unbuf <= my_rom(669);
      when "001010011110" => q_unbuf <= my_rom(670);
      when "001010011111" => q_unbuf <= my_rom(671);
      when "001010100000" => q_unbuf <= my_rom(672);
      when "001010100001" => q_unbuf <= my_rom(673);
      when "001010100010" => q_unbuf <= my_rom(674);
      when "001010100011" => q_unbuf <= my_rom(675);
      when "001010100100" => q_unbuf <= my_rom(676);
      when "001010100101" => q_unbuf <= my_rom(677);
      when "001010100110" => q_unbuf <= my_rom(678);
      when "001010100111" => q_unbuf <= my_rom(679);
      when "001010101000" => q_unbuf <= my_rom(680);
      when "001010101001" => q_unbuf <= my_rom(681);
      when "001010101010" => q_unbuf <= my_rom(682);
      when "001010101011" => q_unbuf <= my_rom(683);
      when "001010101100" => q_unbuf <= my_rom(684);
      when "001010101101" => q_unbuf <= my_rom(685);
      when "001010101110" => q_unbuf <= my_rom(686);
      when "001010101111" => q_unbuf <= my_rom(687);
      when "001010110000" => q_unbuf <= my_rom(688);
      when "001010110001" => q_unbuf <= my_rom(689);
      when "001010110010" => q_unbuf <= my_rom(690);
      when "001010110011" => q_unbuf <= my_rom(691);
      when "001010110100" => q_unbuf <= my_rom(692);
      when "001010110101" => q_unbuf <= my_rom(693);
      when "001010110110" => q_unbuf <= my_rom(694);
      when "001010110111" => q_unbuf <= my_rom(695);
      when "001010111000" => q_unbuf <= my_rom(696);
      when "001010111001" => q_unbuf <= my_rom(697);
      when "001010111010" => q_unbuf <= my_rom(698);
      when "001010111011" => q_unbuf <= my_rom(699);
      when "001010111100" => q_unbuf <= my_rom(700);
      when "001010111101" => q_unbuf <= my_rom(701);
      when "001010111110" => q_unbuf <= my_rom(702);
      when "001010111111" => q_unbuf <= my_rom(703);
      when "001011000000" => q_unbuf <= my_rom(704);
      when "001011000001" => q_unbuf <= my_rom(705);
      when "001011000010" => q_unbuf <= my_rom(706);
      when "001011000011" => q_unbuf <= my_rom(707);
      when "001011000100" => q_unbuf <= my_rom(708);
      when "001011000101" => q_unbuf <= my_rom(709);
      when "001011000110" => q_unbuf <= my_rom(710);
      when "001011000111" => q_unbuf <= my_rom(711);
      when "001011001000" => q_unbuf <= my_rom(712);
      when "001011001001" => q_unbuf <= my_rom(713);
      when "001011001010" => q_unbuf <= my_rom(714);
      when "001011001011" => q_unbuf <= my_rom(715);
      when "001011001100" => q_unbuf <= my_rom(716);
      when "001011001101" => q_unbuf <= my_rom(717);
      when "001011001110" => q_unbuf <= my_rom(718);
      when "001011001111" => q_unbuf <= my_rom(719);
      when "001011010000" => q_unbuf <= my_rom(720);
      when "001011010001" => q_unbuf <= my_rom(721);
      when "001011010010" => q_unbuf <= my_rom(722);
      when "001011010011" => q_unbuf <= my_rom(723);
      when "001011010100" => q_unbuf <= my_rom(724);
      when "001011010101" => q_unbuf <= my_rom(725);
      when "001011010110" => q_unbuf <= my_rom(726);
      when "001011010111" => q_unbuf <= my_rom(727);
      when "001011011000" => q_unbuf <= my_rom(728);
      when "001011011001" => q_unbuf <= my_rom(729);
      when "001011011010" => q_unbuf <= my_rom(730);
      when "001011011011" => q_unbuf <= my_rom(731);
      when "001011011100" => q_unbuf <= my_rom(732);
      when "001011011101" => q_unbuf <= my_rom(733);
      when "001011011110" => q_unbuf <= my_rom(734);
      when "001011011111" => q_unbuf <= my_rom(735);
      when "001011100000" => q_unbuf <= my_rom(736);
      when "001011100001" => q_unbuf <= my_rom(737);
      when "001011100010" => q_unbuf <= my_rom(738);
      when "001011100011" => q_unbuf <= my_rom(739);
      when "001011100100" => q_unbuf <= my_rom(740);
      when "001011100101" => q_unbuf <= my_rom(741);
      when "001011100110" => q_unbuf <= my_rom(742);
      when "001011100111" => q_unbuf <= my_rom(743);
      when "001011101000" => q_unbuf <= my_rom(744);
      when "001011101001" => q_unbuf <= my_rom(745);
      when "001011101010" => q_unbuf <= my_rom(746);
      when "001011101011" => q_unbuf <= my_rom(747);
      when "001011101100" => q_unbuf <= my_rom(748);
      when "001011101101" => q_unbuf <= my_rom(749);
      when "001011101110" => q_unbuf <= my_rom(750);
      when "001011101111" => q_unbuf <= my_rom(751);
      when "001011110000" => q_unbuf <= my_rom(752);
      when "001011110001" => q_unbuf <= my_rom(753);
      when "001011110010" => q_unbuf <= my_rom(754);
      when "001011110011" => q_unbuf <= my_rom(755);
      when "001011110100" => q_unbuf <= my_rom(756);
      when "001011110101" => q_unbuf <= my_rom(757);
      when "001011110110" => q_unbuf <= my_rom(758);
      when "001011110111" => q_unbuf <= my_rom(759);
      when "001011111000" => q_unbuf <= my_rom(760);
      when "001011111001" => q_unbuf <= my_rom(761);
      when "001011111010" => q_unbuf <= my_rom(762);
      when "001011111011" => q_unbuf <= my_rom(763);
      when "001011111100" => q_unbuf <= my_rom(764);
      when "001011111101" => q_unbuf <= my_rom(765);
      when "001011111110" => q_unbuf <= my_rom(766);
      when "001011111111" => q_unbuf <= my_rom(767);
      when "001100000000" => q_unbuf <= my_rom(768);
      when "001100000001" => q_unbuf <= my_rom(769);
      when "001100000010" => q_unbuf <= my_rom(770);
      when "001100000011" => q_unbuf <= my_rom(771);
      when "001100000100" => q_unbuf <= my_rom(772);
      when "001100000101" => q_unbuf <= my_rom(773);
      when "001100000110" => q_unbuf <= my_rom(774);
      when "001100000111" => q_unbuf <= my_rom(775);
      when "001100001000" => q_unbuf <= my_rom(776);
      when "001100001001" => q_unbuf <= my_rom(777);
      when "001100001010" => q_unbuf <= my_rom(778);
      when "001100001011" => q_unbuf <= my_rom(779);
      when "001100001100" => q_unbuf <= my_rom(780);
      when "001100001101" => q_unbuf <= my_rom(781);
      when "001100001110" => q_unbuf <= my_rom(782);
      when "001100001111" => q_unbuf <= my_rom(783);
      when "001100010000" => q_unbuf <= my_rom(784);
      when "001100010001" => q_unbuf <= my_rom(785);
      when "001100010010" => q_unbuf <= my_rom(786);
      when "001100010011" => q_unbuf <= my_rom(787);
      when "001100010100" => q_unbuf <= my_rom(788);
      when "001100010101" => q_unbuf <= my_rom(789);
      when "001100010110" => q_unbuf <= my_rom(790);
      when "001100010111" => q_unbuf <= my_rom(791);
      when "001100011000" => q_unbuf <= my_rom(792);
      when "001100011001" => q_unbuf <= my_rom(793);
      when "001100011010" => q_unbuf <= my_rom(794);
      when "001100011011" => q_unbuf <= my_rom(795);
      when "001100011100" => q_unbuf <= my_rom(796);
      when "001100011101" => q_unbuf <= my_rom(797);
      when "001100011110" => q_unbuf <= my_rom(798);
      when "001100011111" => q_unbuf <= my_rom(799);
      when "001100100000" => q_unbuf <= my_rom(800);
      when "001100100001" => q_unbuf <= my_rom(801);
      when "001100100010" => q_unbuf <= my_rom(802);
      when "001100100011" => q_unbuf <= my_rom(803);
      when "001100100100" => q_unbuf <= my_rom(804);
      when "001100100101" => q_unbuf <= my_rom(805);
      when "001100100110" => q_unbuf <= my_rom(806);
      when "001100100111" => q_unbuf <= my_rom(807);
      when "001100101000" => q_unbuf <= my_rom(808);
      when "001100101001" => q_unbuf <= my_rom(809);
      when "001100101010" => q_unbuf <= my_rom(810);
      when "001100101011" => q_unbuf <= my_rom(811);
      when "001100101100" => q_unbuf <= my_rom(812);
      when "001100101101" => q_unbuf <= my_rom(813);
      when "001100101110" => q_unbuf <= my_rom(814);
      when "001100101111" => q_unbuf <= my_rom(815);
      when "001100110000" => q_unbuf <= my_rom(816);
      when "001100110001" => q_unbuf <= my_rom(817);
      when "001100110010" => q_unbuf <= my_rom(818);
      when "001100110011" => q_unbuf <= my_rom(819);
      when "001100110100" => q_unbuf <= my_rom(820);
      when "001100110101" => q_unbuf <= my_rom(821);
      when "001100110110" => q_unbuf <= my_rom(822);
      when "001100110111" => q_unbuf <= my_rom(823);
      when "001100111000" => q_unbuf <= my_rom(824);
      when "001100111001" => q_unbuf <= my_rom(825);
      when "001100111010" => q_unbuf <= my_rom(826);
      when "001100111011" => q_unbuf <= my_rom(827);
      when "001100111100" => q_unbuf <= my_rom(828);
      when "001100111101" => q_unbuf <= my_rom(829);
      when "001100111110" => q_unbuf <= my_rom(830);
      when "001100111111" => q_unbuf <= my_rom(831);
      when "001101000000" => q_unbuf <= my_rom(832);
      when "001101000001" => q_unbuf <= my_rom(833);
      when "001101000010" => q_unbuf <= my_rom(834);
      when "001101000011" => q_unbuf <= my_rom(835);
      when "001101000100" => q_unbuf <= my_rom(836);
      when "001101000101" => q_unbuf <= my_rom(837);
      when "001101000110" => q_unbuf <= my_rom(838);
      when "001101000111" => q_unbuf <= my_rom(839);
      when "001101001000" => q_unbuf <= my_rom(840);
      when "001101001001" => q_unbuf <= my_rom(841);
      when "001101001010" => q_unbuf <= my_rom(842);
      when "001101001011" => q_unbuf <= my_rom(843);
      when "001101001100" => q_unbuf <= my_rom(844);
      when "001101001101" => q_unbuf <= my_rom(845);
      when "001101001110" => q_unbuf <= my_rom(846);
      when "001101001111" => q_unbuf <= my_rom(847);
      when "001101010000" => q_unbuf <= my_rom(848);
      when "001101010001" => q_unbuf <= my_rom(849);
      when "001101010010" => q_unbuf <= my_rom(850);
      when "001101010011" => q_unbuf <= my_rom(851);
      when "001101010100" => q_unbuf <= my_rom(852);
      when "001101010101" => q_unbuf <= my_rom(853);
      when "001101010110" => q_unbuf <= my_rom(854);
      when "001101010111" => q_unbuf <= my_rom(855);
      when "001101011000" => q_unbuf <= my_rom(856);
      when "001101011001" => q_unbuf <= my_rom(857);
      when "001101011010" => q_unbuf <= my_rom(858);
      when "001101011011" => q_unbuf <= my_rom(859);
      when "001101011100" => q_unbuf <= my_rom(860);
      when "001101011101" => q_unbuf <= my_rom(861);
      when "001101011110" => q_unbuf <= my_rom(862);
      when "001101011111" => q_unbuf <= my_rom(863);
      when "001101100000" => q_unbuf <= my_rom(864);
      when "001101100001" => q_unbuf <= my_rom(865);
      when "001101100010" => q_unbuf <= my_rom(866);
      when "001101100011" => q_unbuf <= my_rom(867);
      when "001101100100" => q_unbuf <= my_rom(868);
      when "001101100101" => q_unbuf <= my_rom(869);
      when "001101100110" => q_unbuf <= my_rom(870);
      when "001101100111" => q_unbuf <= my_rom(871);
      when "001101101000" => q_unbuf <= my_rom(872);
      when "001101101001" => q_unbuf <= my_rom(873);
      when "001101101010" => q_unbuf <= my_rom(874);
      when "001101101011" => q_unbuf <= my_rom(875);
      when "001101101100" => q_unbuf <= my_rom(876);
      when "001101101101" => q_unbuf <= my_rom(877);
      when "001101101110" => q_unbuf <= my_rom(878);
      when "001101101111" => q_unbuf <= my_rom(879);
      when "001101110000" => q_unbuf <= my_rom(880);
      when "001101110001" => q_unbuf <= my_rom(881);
      when "001101110010" => q_unbuf <= my_rom(882);
      when "001101110011" => q_unbuf <= my_rom(883);
      when "001101110100" => q_unbuf <= my_rom(884);
      when "001101110101" => q_unbuf <= my_rom(885);
      when "001101110110" => q_unbuf <= my_rom(886);
      when "001101110111" => q_unbuf <= my_rom(887);
      when "001101111000" => q_unbuf <= my_rom(888);
      when "001101111001" => q_unbuf <= my_rom(889);
      when "001101111010" => q_unbuf <= my_rom(890);
      when "001101111011" => q_unbuf <= my_rom(891);
      when "001101111100" => q_unbuf <= my_rom(892);
      when "001101111101" => q_unbuf <= my_rom(893);
      when "001101111110" => q_unbuf <= my_rom(894);
      when "001101111111" => q_unbuf <= my_rom(895);
      when "001110000000" => q_unbuf <= my_rom(896);
      when "001110000001" => q_unbuf <= my_rom(897);
      when "001110000010" => q_unbuf <= my_rom(898);
      when "001110000011" => q_unbuf <= my_rom(899);
      when "001110000100" => q_unbuf <= my_rom(900);
      when "001110000101" => q_unbuf <= my_rom(901);
      when "001110000110" => q_unbuf <= my_rom(902);
      when "001110000111" => q_unbuf <= my_rom(903);
      when "001110001000" => q_unbuf <= my_rom(904);
      when "001110001001" => q_unbuf <= my_rom(905);
      when "001110001010" => q_unbuf <= my_rom(906);
      when "001110001011" => q_unbuf <= my_rom(907);
      when "001110001100" => q_unbuf <= my_rom(908);
      when "001110001101" => q_unbuf <= my_rom(909);
      when "001110001110" => q_unbuf <= my_rom(910);
      when "001110001111" => q_unbuf <= my_rom(911);
      when "001110010000" => q_unbuf <= my_rom(912);
      when "001110010001" => q_unbuf <= my_rom(913);
      when "001110010010" => q_unbuf <= my_rom(914);
      when "001110010011" => q_unbuf <= my_rom(915);
      when "001110010100" => q_unbuf <= my_rom(916);
      when "001110010101" => q_unbuf <= my_rom(917);
      when "001110010110" => q_unbuf <= my_rom(918);
      when "001110010111" => q_unbuf <= my_rom(919);
      when "001110011000" => q_unbuf <= my_rom(920);
      when "001110011001" => q_unbuf <= my_rom(921);
      when "001110011010" => q_unbuf <= my_rom(922);
      when "001110011011" => q_unbuf <= my_rom(923);
      when "001110011100" => q_unbuf <= my_rom(924);
      when "001110011101" => q_unbuf <= my_rom(925);
      when "001110011110" => q_unbuf <= my_rom(926);
      when "001110011111" => q_unbuf <= my_rom(927);
      when "001110100000" => q_unbuf <= my_rom(928);
      when "001110100001" => q_unbuf <= my_rom(929);
      when "001110100010" => q_unbuf <= my_rom(930);
      when "001110100011" => q_unbuf <= my_rom(931);
      when "001110100100" => q_unbuf <= my_rom(932);
      when "001110100101" => q_unbuf <= my_rom(933);
      when "001110100110" => q_unbuf <= my_rom(934);
      when "001110100111" => q_unbuf <= my_rom(935);
      when "001110101000" => q_unbuf <= my_rom(936);
      when "001110101001" => q_unbuf <= my_rom(937);
      when "001110101010" => q_unbuf <= my_rom(938);
      when "001110101011" => q_unbuf <= my_rom(939);
      when "001110101100" => q_unbuf <= my_rom(940);
      when "001110101101" => q_unbuf <= my_rom(941);
      when "001110101110" => q_unbuf <= my_rom(942);
      when "001110101111" => q_unbuf <= my_rom(943);
      when "001110110000" => q_unbuf <= my_rom(944);
      when "001110110001" => q_unbuf <= my_rom(945);
      when "001110110010" => q_unbuf <= my_rom(946);
      when "001110110011" => q_unbuf <= my_rom(947);
      when "001110110100" => q_unbuf <= my_rom(948);
      when "001110110101" => q_unbuf <= my_rom(949);
      when "001110110110" => q_unbuf <= my_rom(950);
      when "001110110111" => q_unbuf <= my_rom(951);
      when "001110111000" => q_unbuf <= my_rom(952);
      when "001110111001" => q_unbuf <= my_rom(953);
      when "001110111010" => q_unbuf <= my_rom(954);
      when "001110111011" => q_unbuf <= my_rom(955);
      when "001110111100" => q_unbuf <= my_rom(956);
      when "001110111101" => q_unbuf <= my_rom(957);
      when "001110111110" => q_unbuf <= my_rom(958);
      when "001110111111" => q_unbuf <= my_rom(959);
      when "001111000000" => q_unbuf <= my_rom(960);
      when "001111000001" => q_unbuf <= my_rom(961);
      when "001111000010" => q_unbuf <= my_rom(962);
      when "001111000011" => q_unbuf <= my_rom(963);
      when "001111000100" => q_unbuf <= my_rom(964);
      when "001111000101" => q_unbuf <= my_rom(965);
      when "001111000110" => q_unbuf <= my_rom(966);
      when "001111000111" => q_unbuf <= my_rom(967);
      when "001111001000" => q_unbuf <= my_rom(968);
      when "001111001001" => q_unbuf <= my_rom(969);
      when "001111001010" => q_unbuf <= my_rom(970);
      when "001111001011" => q_unbuf <= my_rom(971);
      when "001111001100" => q_unbuf <= my_rom(972);
      when "001111001101" => q_unbuf <= my_rom(973);
      when "001111001110" => q_unbuf <= my_rom(974);
      when "001111001111" => q_unbuf <= my_rom(975);
      when "001111010000" => q_unbuf <= my_rom(976);
      when "001111010001" => q_unbuf <= my_rom(977);
      when "001111010010" => q_unbuf <= my_rom(978);
      when "001111010011" => q_unbuf <= my_rom(979);
      when "001111010100" => q_unbuf <= my_rom(980);
      when "001111010101" => q_unbuf <= my_rom(981);
      when "001111010110" => q_unbuf <= my_rom(982);
      when "001111010111" => q_unbuf <= my_rom(983);
      when "001111011000" => q_unbuf <= my_rom(984);
      when "001111011001" => q_unbuf <= my_rom(985);
      when "001111011010" => q_unbuf <= my_rom(986);
      when "001111011011" => q_unbuf <= my_rom(987);
      when "001111011100" => q_unbuf <= my_rom(988);
      when "001111011101" => q_unbuf <= my_rom(989);
      when "001111011110" => q_unbuf <= my_rom(990);
      when "001111011111" => q_unbuf <= my_rom(991);
      when "001111100000" => q_unbuf <= my_rom(992);
      when "001111100001" => q_unbuf <= my_rom(993);
      when "001111100010" => q_unbuf <= my_rom(994);
      when "001111100011" => q_unbuf <= my_rom(995);
      when "001111100100" => q_unbuf <= my_rom(996);
      when "001111100101" => q_unbuf <= my_rom(997);
      when "001111100110" => q_unbuf <= my_rom(998);
      when "001111100111" => q_unbuf <= my_rom(999);
      when "001111101000" => q_unbuf <= my_rom(1000);
      when "001111101001" => q_unbuf <= my_rom(1001);
      when "001111101010" => q_unbuf <= my_rom(1002);
      when "001111101011" => q_unbuf <= my_rom(1003);
      when "001111101100" => q_unbuf <= my_rom(1004);
      when "001111101101" => q_unbuf <= my_rom(1005);
      when "001111101110" => q_unbuf <= my_rom(1006);
      when "001111101111" => q_unbuf <= my_rom(1007);
      when "001111110000" => q_unbuf <= my_rom(1008);
      when "001111110001" => q_unbuf <= my_rom(1009);
      when "001111110010" => q_unbuf <= my_rom(1010);
      when "001111110011" => q_unbuf <= my_rom(1011);
      when "001111110100" => q_unbuf <= my_rom(1012);
      when "001111110101" => q_unbuf <= my_rom(1013);
      when "001111110110" => q_unbuf <= my_rom(1014);
      when "001111110111" => q_unbuf <= my_rom(1015);
      when "001111111000" => q_unbuf <= my_rom(1016);
      when "001111111001" => q_unbuf <= my_rom(1017);
      when "001111111010" => q_unbuf <= my_rom(1018);
      when "001111111011" => q_unbuf <= my_rom(1019);
      when "001111111100" => q_unbuf <= my_rom(1020);
      when "001111111101" => q_unbuf <= my_rom(1021);
      when "001111111110" => q_unbuf <= my_rom(1022);
      when "001111111111" => q_unbuf <= my_rom(1023);
      when "010000000000" => q_unbuf <= my_rom(1024);
      when "010000000001" => q_unbuf <= my_rom(1025);
      when "010000000010" => q_unbuf <= my_rom(1026);
      when "010000000011" => q_unbuf <= my_rom(1027);
      when "010000000100" => q_unbuf <= my_rom(1028);
      when "010000000101" => q_unbuf <= my_rom(1029);
      when "010000000110" => q_unbuf <= my_rom(1030);
      when "010000000111" => q_unbuf <= my_rom(1031);
      when "010000001000" => q_unbuf <= my_rom(1032);
      when "010000001001" => q_unbuf <= my_rom(1033);
      when "010000001010" => q_unbuf <= my_rom(1034);
      when "010000001011" => q_unbuf <= my_rom(1035);
      when "010000001100" => q_unbuf <= my_rom(1036);
      when "010000001101" => q_unbuf <= my_rom(1037);
      when "010000001110" => q_unbuf <= my_rom(1038);
      when "010000001111" => q_unbuf <= my_rom(1039);
      when "010000010000" => q_unbuf <= my_rom(1040);
      when "010000010001" => q_unbuf <= my_rom(1041);
      when "010000010010" => q_unbuf <= my_rom(1042);
      when "010000010011" => q_unbuf <= my_rom(1043);
      when "010000010100" => q_unbuf <= my_rom(1044);
      when "010000010101" => q_unbuf <= my_rom(1045);
      when "010000010110" => q_unbuf <= my_rom(1046);
      when "010000010111" => q_unbuf <= my_rom(1047);
      when "010000011000" => q_unbuf <= my_rom(1048);
      when "010000011001" => q_unbuf <= my_rom(1049);
      when "010000011010" => q_unbuf <= my_rom(1050);
      when "010000011011" => q_unbuf <= my_rom(1051);
      when "010000011100" => q_unbuf <= my_rom(1052);
      when "010000011101" => q_unbuf <= my_rom(1053);
      when "010000011110" => q_unbuf <= my_rom(1054);
      when "010000011111" => q_unbuf <= my_rom(1055);
      when "010000100000" => q_unbuf <= my_rom(1056);
      when "010000100001" => q_unbuf <= my_rom(1057);
      when "010000100010" => q_unbuf <= my_rom(1058);
      when "010000100011" => q_unbuf <= my_rom(1059);
      when "010000100100" => q_unbuf <= my_rom(1060);
      when "010000100101" => q_unbuf <= my_rom(1061);
      when "010000100110" => q_unbuf <= my_rom(1062);
      when "010000100111" => q_unbuf <= my_rom(1063);
      when "010000101000" => q_unbuf <= my_rom(1064);
      when "010000101001" => q_unbuf <= my_rom(1065);
      when "010000101010" => q_unbuf <= my_rom(1066);
      when "010000101011" => q_unbuf <= my_rom(1067);
      when "010000101100" => q_unbuf <= my_rom(1068);
      when "010000101101" => q_unbuf <= my_rom(1069);
      when "010000101110" => q_unbuf <= my_rom(1070);
      when "010000101111" => q_unbuf <= my_rom(1071);
      when "010000110000" => q_unbuf <= my_rom(1072);
      when "010000110001" => q_unbuf <= my_rom(1073);
      when "010000110010" => q_unbuf <= my_rom(1074);
      when "010000110011" => q_unbuf <= my_rom(1075);
      when "010000110100" => q_unbuf <= my_rom(1076);
      when "010000110101" => q_unbuf <= my_rom(1077);
      when "010000110110" => q_unbuf <= my_rom(1078);
      when "010000110111" => q_unbuf <= my_rom(1079);
      when "010000111000" => q_unbuf <= my_rom(1080);
      when "010000111001" => q_unbuf <= my_rom(1081);
      when "010000111010" => q_unbuf <= my_rom(1082);
      when "010000111011" => q_unbuf <= my_rom(1083);
      when "010000111100" => q_unbuf <= my_rom(1084);
      when "010000111101" => q_unbuf <= my_rom(1085);
      when "010000111110" => q_unbuf <= my_rom(1086);
      when "010000111111" => q_unbuf <= my_rom(1087);
      when "010001000000" => q_unbuf <= my_rom(1088);
      when "010001000001" => q_unbuf <= my_rom(1089);
      when "010001000010" => q_unbuf <= my_rom(1090);
      when "010001000011" => q_unbuf <= my_rom(1091);
      when "010001000100" => q_unbuf <= my_rom(1092);
      when "010001000101" => q_unbuf <= my_rom(1093);
      when "010001000110" => q_unbuf <= my_rom(1094);
      when "010001000111" => q_unbuf <= my_rom(1095);
      when "010001001000" => q_unbuf <= my_rom(1096);
      when "010001001001" => q_unbuf <= my_rom(1097);
      when "010001001010" => q_unbuf <= my_rom(1098);
      when "010001001011" => q_unbuf <= my_rom(1099);
      when "010001001100" => q_unbuf <= my_rom(1100);
      when "010001001101" => q_unbuf <= my_rom(1101);
      when "010001001110" => q_unbuf <= my_rom(1102);
      when "010001001111" => q_unbuf <= my_rom(1103);
      when "010001010000" => q_unbuf <= my_rom(1104);
      when "010001010001" => q_unbuf <= my_rom(1105);
      when "010001010010" => q_unbuf <= my_rom(1106);
      when "010001010011" => q_unbuf <= my_rom(1107);
      when "010001010100" => q_unbuf <= my_rom(1108);
      when "010001010101" => q_unbuf <= my_rom(1109);
      when "010001010110" => q_unbuf <= my_rom(1110);
      when "010001010111" => q_unbuf <= my_rom(1111);
      when "010001011000" => q_unbuf <= my_rom(1112);
      when "010001011001" => q_unbuf <= my_rom(1113);
      when "010001011010" => q_unbuf <= my_rom(1114);
      when "010001011011" => q_unbuf <= my_rom(1115);
      when "010001011100" => q_unbuf <= my_rom(1116);
      when "010001011101" => q_unbuf <= my_rom(1117);
      when "010001011110" => q_unbuf <= my_rom(1118);
      when "010001011111" => q_unbuf <= my_rom(1119);
      when "010001100000" => q_unbuf <= my_rom(1120);
      when "010001100001" => q_unbuf <= my_rom(1121);
      when "010001100010" => q_unbuf <= my_rom(1122);
      when "010001100011" => q_unbuf <= my_rom(1123);
      when "010001100100" => q_unbuf <= my_rom(1124);
      when "010001100101" => q_unbuf <= my_rom(1125);
      when "010001100110" => q_unbuf <= my_rom(1126);
      when "010001100111" => q_unbuf <= my_rom(1127);
      when "010001101000" => q_unbuf <= my_rom(1128);
      when "010001101001" => q_unbuf <= my_rom(1129);
      when "010001101010" => q_unbuf <= my_rom(1130);
      when "010001101011" => q_unbuf <= my_rom(1131);
      when "010001101100" => q_unbuf <= my_rom(1132);
      when "010001101101" => q_unbuf <= my_rom(1133);
      when "010001101110" => q_unbuf <= my_rom(1134);
      when "010001101111" => q_unbuf <= my_rom(1135);
      when "010001110000" => q_unbuf <= my_rom(1136);
      when "010001110001" => q_unbuf <= my_rom(1137);
      when "010001110010" => q_unbuf <= my_rom(1138);
      when "010001110011" => q_unbuf <= my_rom(1139);
      when "010001110100" => q_unbuf <= my_rom(1140);
      when "010001110101" => q_unbuf <= my_rom(1141);
      when "010001110110" => q_unbuf <= my_rom(1142);
      when "010001110111" => q_unbuf <= my_rom(1143);
      when "010001111000" => q_unbuf <= my_rom(1144);
      when "010001111001" => q_unbuf <= my_rom(1145);
      when "010001111010" => q_unbuf <= my_rom(1146);
      when "010001111011" => q_unbuf <= my_rom(1147);
      when "010001111100" => q_unbuf <= my_rom(1148);
      when "010001111101" => q_unbuf <= my_rom(1149);
      when "010001111110" => q_unbuf <= my_rom(1150);
      when "010001111111" => q_unbuf <= my_rom(1151);
      when "010010000000" => q_unbuf <= my_rom(1152);
      when "010010000001" => q_unbuf <= my_rom(1153);
      when "010010000010" => q_unbuf <= my_rom(1154);
      when "010010000011" => q_unbuf <= my_rom(1155);
      when "010010000100" => q_unbuf <= my_rom(1156);
      when "010010000101" => q_unbuf <= my_rom(1157);
      when "010010000110" => q_unbuf <= my_rom(1158);
      when "010010000111" => q_unbuf <= my_rom(1159);
      when "010010001000" => q_unbuf <= my_rom(1160);
      when "010010001001" => q_unbuf <= my_rom(1161);
      when "010010001010" => q_unbuf <= my_rom(1162);
      when "010010001011" => q_unbuf <= my_rom(1163);
      when "010010001100" => q_unbuf <= my_rom(1164);
      when "010010001101" => q_unbuf <= my_rom(1165);
      when "010010001110" => q_unbuf <= my_rom(1166);
      when "010010001111" => q_unbuf <= my_rom(1167);
      when "010010010000" => q_unbuf <= my_rom(1168);
      when "010010010001" => q_unbuf <= my_rom(1169);
      when "010010010010" => q_unbuf <= my_rom(1170);
      when "010010010011" => q_unbuf <= my_rom(1171);
      when "010010010100" => q_unbuf <= my_rom(1172);
      when "010010010101" => q_unbuf <= my_rom(1173);
      when "010010010110" => q_unbuf <= my_rom(1174);
      when "010010010111" => q_unbuf <= my_rom(1175);
      when "010010011000" => q_unbuf <= my_rom(1176);
      when "010010011001" => q_unbuf <= my_rom(1177);
      when "010010011010" => q_unbuf <= my_rom(1178);
      when "010010011011" => q_unbuf <= my_rom(1179);
      when "010010011100" => q_unbuf <= my_rom(1180);
      when "010010011101" => q_unbuf <= my_rom(1181);
      when "010010011110" => q_unbuf <= my_rom(1182);
      when "010010011111" => q_unbuf <= my_rom(1183);
      when "010010100000" => q_unbuf <= my_rom(1184);
      when "010010100001" => q_unbuf <= my_rom(1185);
      when "010010100010" => q_unbuf <= my_rom(1186);
      when "010010100011" => q_unbuf <= my_rom(1187);
      when "010010100100" => q_unbuf <= my_rom(1188);
      when "010010100101" => q_unbuf <= my_rom(1189);
      when "010010100110" => q_unbuf <= my_rom(1190);
      when "010010100111" => q_unbuf <= my_rom(1191);
      when "010010101000" => q_unbuf <= my_rom(1192);
      when "010010101001" => q_unbuf <= my_rom(1193);
      when "010010101010" => q_unbuf <= my_rom(1194);
      when "010010101011" => q_unbuf <= my_rom(1195);
      when "010010101100" => q_unbuf <= my_rom(1196);
      when "010010101101" => q_unbuf <= my_rom(1197);
      when "010010101110" => q_unbuf <= my_rom(1198);
      when "010010101111" => q_unbuf <= my_rom(1199);
      when "010010110000" => q_unbuf <= my_rom(1200);
      when "010010110001" => q_unbuf <= my_rom(1201);
      when "010010110010" => q_unbuf <= my_rom(1202);
      when "010010110011" => q_unbuf <= my_rom(1203);
      when "010010110100" => q_unbuf <= my_rom(1204);
      when "010010110101" => q_unbuf <= my_rom(1205);
      when "010010110110" => q_unbuf <= my_rom(1206);
      when "010010110111" => q_unbuf <= my_rom(1207);
      when "010010111000" => q_unbuf <= my_rom(1208);
      when "010010111001" => q_unbuf <= my_rom(1209);
      when "010010111010" => q_unbuf <= my_rom(1210);
      when "010010111011" => q_unbuf <= my_rom(1211);
      when "010010111100" => q_unbuf <= my_rom(1212);
      when "010010111101" => q_unbuf <= my_rom(1213);
      when "010010111110" => q_unbuf <= my_rom(1214);
      when "010010111111" => q_unbuf <= my_rom(1215);
      when "010011000000" => q_unbuf <= my_rom(1216);
      when "010011000001" => q_unbuf <= my_rom(1217);
      when "010011000010" => q_unbuf <= my_rom(1218);
      when "010011000011" => q_unbuf <= my_rom(1219);
      when "010011000100" => q_unbuf <= my_rom(1220);
      when "010011000101" => q_unbuf <= my_rom(1221);
      when "010011000110" => q_unbuf <= my_rom(1222);
      when "010011000111" => q_unbuf <= my_rom(1223);
      when "010011001000" => q_unbuf <= my_rom(1224);
      when "010011001001" => q_unbuf <= my_rom(1225);
      when "010011001010" => q_unbuf <= my_rom(1226);
      when "010011001011" => q_unbuf <= my_rom(1227);
      when "010011001100" => q_unbuf <= my_rom(1228);
      when "010011001101" => q_unbuf <= my_rom(1229);
      when "010011001110" => q_unbuf <= my_rom(1230);
      when "010011001111" => q_unbuf <= my_rom(1231);
      when "010011010000" => q_unbuf <= my_rom(1232);
      when "010011010001" => q_unbuf <= my_rom(1233);
      when "010011010010" => q_unbuf <= my_rom(1234);
      when "010011010011" => q_unbuf <= my_rom(1235);
      when "010011010100" => q_unbuf <= my_rom(1236);
      when "010011010101" => q_unbuf <= my_rom(1237);
      when "010011010110" => q_unbuf <= my_rom(1238);
      when "010011010111" => q_unbuf <= my_rom(1239);
      when "010011011000" => q_unbuf <= my_rom(1240);
      when "010011011001" => q_unbuf <= my_rom(1241);
      when "010011011010" => q_unbuf <= my_rom(1242);
      when "010011011011" => q_unbuf <= my_rom(1243);
      when "010011011100" => q_unbuf <= my_rom(1244);
      when "010011011101" => q_unbuf <= my_rom(1245);
      when "010011011110" => q_unbuf <= my_rom(1246);
      when "010011011111" => q_unbuf <= my_rom(1247);
      when "010011100000" => q_unbuf <= my_rom(1248);
      when "010011100001" => q_unbuf <= my_rom(1249);
      when "010011100010" => q_unbuf <= my_rom(1250);
      when "010011100011" => q_unbuf <= my_rom(1251);
      when "010011100100" => q_unbuf <= my_rom(1252);
      when "010011100101" => q_unbuf <= my_rom(1253);
      when "010011100110" => q_unbuf <= my_rom(1254);
      when "010011100111" => q_unbuf <= my_rom(1255);
      when "010011101000" => q_unbuf <= my_rom(1256);
      when "010011101001" => q_unbuf <= my_rom(1257);
      when "010011101010" => q_unbuf <= my_rom(1258);
      when "010011101011" => q_unbuf <= my_rom(1259);
      when "010011101100" => q_unbuf <= my_rom(1260);
      when "010011101101" => q_unbuf <= my_rom(1261);
      when "010011101110" => q_unbuf <= my_rom(1262);
      when "010011101111" => q_unbuf <= my_rom(1263);
      when "010011110000" => q_unbuf <= my_rom(1264);
      when "010011110001" => q_unbuf <= my_rom(1265);
      when "010011110010" => q_unbuf <= my_rom(1266);
      when "010011110011" => q_unbuf <= my_rom(1267);
      when "010011110100" => q_unbuf <= my_rom(1268);
      when "010011110101" => q_unbuf <= my_rom(1269);
      when "010011110110" => q_unbuf <= my_rom(1270);
      when "010011110111" => q_unbuf <= my_rom(1271);
      when "010011111000" => q_unbuf <= my_rom(1272);
      when "010011111001" => q_unbuf <= my_rom(1273);
      when "010011111010" => q_unbuf <= my_rom(1274);
      when "010011111011" => q_unbuf <= my_rom(1275);
      when "010011111100" => q_unbuf <= my_rom(1276);
      when "010011111101" => q_unbuf <= my_rom(1277);
      when "010011111110" => q_unbuf <= my_rom(1278);
      when "010011111111" => q_unbuf <= my_rom(1279);
      when "010100000000" => q_unbuf <= my_rom(1280);
      when "010100000001" => q_unbuf <= my_rom(1281);
      when "010100000010" => q_unbuf <= my_rom(1282);
      when "010100000011" => q_unbuf <= my_rom(1283);
      when "010100000100" => q_unbuf <= my_rom(1284);
      when "010100000101" => q_unbuf <= my_rom(1285);
      when "010100000110" => q_unbuf <= my_rom(1286);
      when "010100000111" => q_unbuf <= my_rom(1287);
      when "010100001000" => q_unbuf <= my_rom(1288);
      when "010100001001" => q_unbuf <= my_rom(1289);
      when "010100001010" => q_unbuf <= my_rom(1290);
      when "010100001011" => q_unbuf <= my_rom(1291);
      when "010100001100" => q_unbuf <= my_rom(1292);
      when "010100001101" => q_unbuf <= my_rom(1293);
      when "010100001110" => q_unbuf <= my_rom(1294);
      when "010100001111" => q_unbuf <= my_rom(1295);
      when "010100010000" => q_unbuf <= my_rom(1296);
      when "010100010001" => q_unbuf <= my_rom(1297);
      when "010100010010" => q_unbuf <= my_rom(1298);
      when "010100010011" => q_unbuf <= my_rom(1299);
      when "010100010100" => q_unbuf <= my_rom(1300);
      when "010100010101" => q_unbuf <= my_rom(1301);
      when "010100010110" => q_unbuf <= my_rom(1302);
      when "010100010111" => q_unbuf <= my_rom(1303);
      when "010100011000" => q_unbuf <= my_rom(1304);
      when "010100011001" => q_unbuf <= my_rom(1305);
      when "010100011010" => q_unbuf <= my_rom(1306);
      when "010100011011" => q_unbuf <= my_rom(1307);
      when "010100011100" => q_unbuf <= my_rom(1308);
      when "010100011101" => q_unbuf <= my_rom(1309);
      when "010100011110" => q_unbuf <= my_rom(1310);
      when "010100011111" => q_unbuf <= my_rom(1311);
      when "010100100000" => q_unbuf <= my_rom(1312);
      when "010100100001" => q_unbuf <= my_rom(1313);
      when "010100100010" => q_unbuf <= my_rom(1314);
      when "010100100011" => q_unbuf <= my_rom(1315);
      when "010100100100" => q_unbuf <= my_rom(1316);
      when "010100100101" => q_unbuf <= my_rom(1317);
      when "010100100110" => q_unbuf <= my_rom(1318);
      when "010100100111" => q_unbuf <= my_rom(1319);
      when "010100101000" => q_unbuf <= my_rom(1320);
      when "010100101001" => q_unbuf <= my_rom(1321);
      when "010100101010" => q_unbuf <= my_rom(1322);
      when "010100101011" => q_unbuf <= my_rom(1323);
      when "010100101100" => q_unbuf <= my_rom(1324);
      when "010100101101" => q_unbuf <= my_rom(1325);
      when "010100101110" => q_unbuf <= my_rom(1326);
      when "010100101111" => q_unbuf <= my_rom(1327);
      when "010100110000" => q_unbuf <= my_rom(1328);
      when "010100110001" => q_unbuf <= my_rom(1329);
      when "010100110010" => q_unbuf <= my_rom(1330);
      when "010100110011" => q_unbuf <= my_rom(1331);
      when "010100110100" => q_unbuf <= my_rom(1332);
      when "010100110101" => q_unbuf <= my_rom(1333);
      when "010100110110" => q_unbuf <= my_rom(1334);
      when "010100110111" => q_unbuf <= my_rom(1335);
      when "010100111000" => q_unbuf <= my_rom(1336);
      when "010100111001" => q_unbuf <= my_rom(1337);
      when "010100111010" => q_unbuf <= my_rom(1338);
      when "010100111011" => q_unbuf <= my_rom(1339);
      when "010100111100" => q_unbuf <= my_rom(1340);
      when "010100111101" => q_unbuf <= my_rom(1341);
      when "010100111110" => q_unbuf <= my_rom(1342);
      when "010100111111" => q_unbuf <= my_rom(1343);
      when "010101000000" => q_unbuf <= my_rom(1344);
      when "010101000001" => q_unbuf <= my_rom(1345);
      when "010101000010" => q_unbuf <= my_rom(1346);
      when "010101000011" => q_unbuf <= my_rom(1347);
      when "010101000100" => q_unbuf <= my_rom(1348);
      when "010101000101" => q_unbuf <= my_rom(1349);
      when "010101000110" => q_unbuf <= my_rom(1350);
      when "010101000111" => q_unbuf <= my_rom(1351);
      when "010101001000" => q_unbuf <= my_rom(1352);
      when "010101001001" => q_unbuf <= my_rom(1353);
      when "010101001010" => q_unbuf <= my_rom(1354);
      when "010101001011" => q_unbuf <= my_rom(1355);
      when "010101001100" => q_unbuf <= my_rom(1356);
      when "010101001101" => q_unbuf <= my_rom(1357);
      when "010101001110" => q_unbuf <= my_rom(1358);
      when "010101001111" => q_unbuf <= my_rom(1359);
      when "010101010000" => q_unbuf <= my_rom(1360);
      when "010101010001" => q_unbuf <= my_rom(1361);
      when "010101010010" => q_unbuf <= my_rom(1362);
      when "010101010011" => q_unbuf <= my_rom(1363);
      when "010101010100" => q_unbuf <= my_rom(1364);
      when "010101010101" => q_unbuf <= my_rom(1365);
      when "010101010110" => q_unbuf <= my_rom(1366);
      when "010101010111" => q_unbuf <= my_rom(1367);
      when "010101011000" => q_unbuf <= my_rom(1368);
      when "010101011001" => q_unbuf <= my_rom(1369);
      when "010101011010" => q_unbuf <= my_rom(1370);
      when "010101011011" => q_unbuf <= my_rom(1371);
      when "010101011100" => q_unbuf <= my_rom(1372);
      when "010101011101" => q_unbuf <= my_rom(1373);
      when "010101011110" => q_unbuf <= my_rom(1374);
      when "010101011111" => q_unbuf <= my_rom(1375);
      when "010101100000" => q_unbuf <= my_rom(1376);
      when "010101100001" => q_unbuf <= my_rom(1377);
      when "010101100010" => q_unbuf <= my_rom(1378);
      when "010101100011" => q_unbuf <= my_rom(1379);
      when "010101100100" => q_unbuf <= my_rom(1380);
      when "010101100101" => q_unbuf <= my_rom(1381);
      when "010101100110" => q_unbuf <= my_rom(1382);
      when "010101100111" => q_unbuf <= my_rom(1383);
      when "010101101000" => q_unbuf <= my_rom(1384);
      when "010101101001" => q_unbuf <= my_rom(1385);
      when "010101101010" => q_unbuf <= my_rom(1386);
      when "010101101011" => q_unbuf <= my_rom(1387);
      when "010101101100" => q_unbuf <= my_rom(1388);
      when "010101101101" => q_unbuf <= my_rom(1389);
      when "010101101110" => q_unbuf <= my_rom(1390);
      when "010101101111" => q_unbuf <= my_rom(1391);
      when "010101110000" => q_unbuf <= my_rom(1392);
      when "010101110001" => q_unbuf <= my_rom(1393);
      when "010101110010" => q_unbuf <= my_rom(1394);
      when "010101110011" => q_unbuf <= my_rom(1395);
      when "010101110100" => q_unbuf <= my_rom(1396);
      when "010101110101" => q_unbuf <= my_rom(1397);
      when "010101110110" => q_unbuf <= my_rom(1398);
      when "010101110111" => q_unbuf <= my_rom(1399);
      when "010101111000" => q_unbuf <= my_rom(1400);
      when "010101111001" => q_unbuf <= my_rom(1401);
      when "010101111010" => q_unbuf <= my_rom(1402);
      when "010101111011" => q_unbuf <= my_rom(1403);
      when "010101111100" => q_unbuf <= my_rom(1404);
      when "010101111101" => q_unbuf <= my_rom(1405);
      when "010101111110" => q_unbuf <= my_rom(1406);
      when "010101111111" => q_unbuf <= my_rom(1407);
      when "010110000000" => q_unbuf <= my_rom(1408);
      when "010110000001" => q_unbuf <= my_rom(1409);
      when "010110000010" => q_unbuf <= my_rom(1410);
      when "010110000011" => q_unbuf <= my_rom(1411);
      when "010110000100" => q_unbuf <= my_rom(1412);
      when "010110000101" => q_unbuf <= my_rom(1413);
      when "010110000110" => q_unbuf <= my_rom(1414);
      when "010110000111" => q_unbuf <= my_rom(1415);
      when "010110001000" => q_unbuf <= my_rom(1416);
      when "010110001001" => q_unbuf <= my_rom(1417);
      when "010110001010" => q_unbuf <= my_rom(1418);
      when "010110001011" => q_unbuf <= my_rom(1419);
      when "010110001100" => q_unbuf <= my_rom(1420);
      when "010110001101" => q_unbuf <= my_rom(1421);
      when "010110001110" => q_unbuf <= my_rom(1422);
      when "010110001111" => q_unbuf <= my_rom(1423);
      when "010110010000" => q_unbuf <= my_rom(1424);
      when "010110010001" => q_unbuf <= my_rom(1425);
      when "010110010010" => q_unbuf <= my_rom(1426);
      when "010110010011" => q_unbuf <= my_rom(1427);
      when "010110010100" => q_unbuf <= my_rom(1428);
      when "010110010101" => q_unbuf <= my_rom(1429);
      when "010110010110" => q_unbuf <= my_rom(1430);
      when "010110010111" => q_unbuf <= my_rom(1431);
      when "010110011000" => q_unbuf <= my_rom(1432);
      when "010110011001" => q_unbuf <= my_rom(1433);
      when "010110011010" => q_unbuf <= my_rom(1434);
      when "010110011011" => q_unbuf <= my_rom(1435);
      when "010110011100" => q_unbuf <= my_rom(1436);
      when "010110011101" => q_unbuf <= my_rom(1437);
      when "010110011110" => q_unbuf <= my_rom(1438);
      when "010110011111" => q_unbuf <= my_rom(1439);
      when "010110100000" => q_unbuf <= my_rom(1440);
      when "010110100001" => q_unbuf <= my_rom(1441);
      when "010110100010" => q_unbuf <= my_rom(1442);
      when "010110100011" => q_unbuf <= my_rom(1443);
      when "010110100100" => q_unbuf <= my_rom(1444);
      when "010110100101" => q_unbuf <= my_rom(1445);
      when "010110100110" => q_unbuf <= my_rom(1446);
      when "010110100111" => q_unbuf <= my_rom(1447);
      when "010110101000" => q_unbuf <= my_rom(1448);
      when "010110101001" => q_unbuf <= my_rom(1449);
      when "010110101010" => q_unbuf <= my_rom(1450);
      when "010110101011" => q_unbuf <= my_rom(1451);
      when "010110101100" => q_unbuf <= my_rom(1452);
      when "010110101101" => q_unbuf <= my_rom(1453);
      when "010110101110" => q_unbuf <= my_rom(1454);
      when "010110101111" => q_unbuf <= my_rom(1455);
      when "010110110000" => q_unbuf <= my_rom(1456);
      when "010110110001" => q_unbuf <= my_rom(1457);
      when "010110110010" => q_unbuf <= my_rom(1458);
      when "010110110011" => q_unbuf <= my_rom(1459);
      when "010110110100" => q_unbuf <= my_rom(1460);
      when "010110110101" => q_unbuf <= my_rom(1461);
      when "010110110110" => q_unbuf <= my_rom(1462);
      when "010110110111" => q_unbuf <= my_rom(1463);
      when "010110111000" => q_unbuf <= my_rom(1464);
      when "010110111001" => q_unbuf <= my_rom(1465);
      when "010110111010" => q_unbuf <= my_rom(1466);
      when "010110111011" => q_unbuf <= my_rom(1467);
      when "010110111100" => q_unbuf <= my_rom(1468);
      when "010110111101" => q_unbuf <= my_rom(1469);
      when "010110111110" => q_unbuf <= my_rom(1470);
      when "010110111111" => q_unbuf <= my_rom(1471);
      when "010111000000" => q_unbuf <= my_rom(1472);
      when "010111000001" => q_unbuf <= my_rom(1473);
      when "010111000010" => q_unbuf <= my_rom(1474);
      when "010111000011" => q_unbuf <= my_rom(1475);
      when "010111000100" => q_unbuf <= my_rom(1476);
      when "010111000101" => q_unbuf <= my_rom(1477);
      when "010111000110" => q_unbuf <= my_rom(1478);
      when "010111000111" => q_unbuf <= my_rom(1479);
      when "010111001000" => q_unbuf <= my_rom(1480);
      when "010111001001" => q_unbuf <= my_rom(1481);
      when "010111001010" => q_unbuf <= my_rom(1482);
      when "010111001011" => q_unbuf <= my_rom(1483);
      when "010111001100" => q_unbuf <= my_rom(1484);
      when "010111001101" => q_unbuf <= my_rom(1485);
      when "010111001110" => q_unbuf <= my_rom(1486);
      when "010111001111" => q_unbuf <= my_rom(1487);
      when "010111010000" => q_unbuf <= my_rom(1488);
      when "010111010001" => q_unbuf <= my_rom(1489);
      when "010111010010" => q_unbuf <= my_rom(1490);
      when "010111010011" => q_unbuf <= my_rom(1491);
      when "010111010100" => q_unbuf <= my_rom(1492);
      when "010111010101" => q_unbuf <= my_rom(1493);
      when "010111010110" => q_unbuf <= my_rom(1494);
      when "010111010111" => q_unbuf <= my_rom(1495);
      when "010111011000" => q_unbuf <= my_rom(1496);
      when "010111011001" => q_unbuf <= my_rom(1497);
      when "010111011010" => q_unbuf <= my_rom(1498);
      when "010111011011" => q_unbuf <= my_rom(1499);
      when "010111011100" => q_unbuf <= my_rom(1500);
      when "010111011101" => q_unbuf <= my_rom(1501);
      when "010111011110" => q_unbuf <= my_rom(1502);
      when "010111011111" => q_unbuf <= my_rom(1503);
      when "010111100000" => q_unbuf <= my_rom(1504);
      when "010111100001" => q_unbuf <= my_rom(1505);
      when "010111100010" => q_unbuf <= my_rom(1506);
      when "010111100011" => q_unbuf <= my_rom(1507);
      when "010111100100" => q_unbuf <= my_rom(1508);
      when "010111100101" => q_unbuf <= my_rom(1509);
      when "010111100110" => q_unbuf <= my_rom(1510);
      when "010111100111" => q_unbuf <= my_rom(1511);
      when "010111101000" => q_unbuf <= my_rom(1512);
      when "010111101001" => q_unbuf <= my_rom(1513);
      when "010111101010" => q_unbuf <= my_rom(1514);
      when "010111101011" => q_unbuf <= my_rom(1515);
      when "010111101100" => q_unbuf <= my_rom(1516);
      when "010111101101" => q_unbuf <= my_rom(1517);
      when "010111101110" => q_unbuf <= my_rom(1518);
      when "010111101111" => q_unbuf <= my_rom(1519);
      when "010111110000" => q_unbuf <= my_rom(1520);
      when "010111110001" => q_unbuf <= my_rom(1521);
      when "010111110010" => q_unbuf <= my_rom(1522);
      when "010111110011" => q_unbuf <= my_rom(1523);
      when "010111110100" => q_unbuf <= my_rom(1524);
      when "010111110101" => q_unbuf <= my_rom(1525);
      when "010111110110" => q_unbuf <= my_rom(1526);
      when "010111110111" => q_unbuf <= my_rom(1527);
      when "010111111000" => q_unbuf <= my_rom(1528);
      when "010111111001" => q_unbuf <= my_rom(1529);
      when "010111111010" => q_unbuf <= my_rom(1530);
      when "010111111011" => q_unbuf <= my_rom(1531);
      when "010111111100" => q_unbuf <= my_rom(1532);
      when "010111111101" => q_unbuf <= my_rom(1533);
      when "010111111110" => q_unbuf <= my_rom(1534);
      when "010111111111" => q_unbuf <= my_rom(1535);
      when "011000000000" => q_unbuf <= my_rom(1536);
      when "011000000001" => q_unbuf <= my_rom(1537);
      when "011000000010" => q_unbuf <= my_rom(1538);
      when "011000000011" => q_unbuf <= my_rom(1539);
      when "011000000100" => q_unbuf <= my_rom(1540);
      when "011000000101" => q_unbuf <= my_rom(1541);
      when "011000000110" => q_unbuf <= my_rom(1542);
      when "011000000111" => q_unbuf <= my_rom(1543);
      when "011000001000" => q_unbuf <= my_rom(1544);
      when "011000001001" => q_unbuf <= my_rom(1545);
      when "011000001010" => q_unbuf <= my_rom(1546);
      when "011000001011" => q_unbuf <= my_rom(1547);
      when "011000001100" => q_unbuf <= my_rom(1548);
      when "011000001101" => q_unbuf <= my_rom(1549);
      when "011000001110" => q_unbuf <= my_rom(1550);
      when "011000001111" => q_unbuf <= my_rom(1551);
      when "011000010000" => q_unbuf <= my_rom(1552);
      when "011000010001" => q_unbuf <= my_rom(1553);
      when "011000010010" => q_unbuf <= my_rom(1554);
      when "011000010011" => q_unbuf <= my_rom(1555);
      when "011000010100" => q_unbuf <= my_rom(1556);
      when "011000010101" => q_unbuf <= my_rom(1557);
      when "011000010110" => q_unbuf <= my_rom(1558);
      when "011000010111" => q_unbuf <= my_rom(1559);
      when "011000011000" => q_unbuf <= my_rom(1560);
      when "011000011001" => q_unbuf <= my_rom(1561);
      when "011000011010" => q_unbuf <= my_rom(1562);
      when "011000011011" => q_unbuf <= my_rom(1563);
      when "011000011100" => q_unbuf <= my_rom(1564);
      when "011000011101" => q_unbuf <= my_rom(1565);
      when "011000011110" => q_unbuf <= my_rom(1566);
      when "011000011111" => q_unbuf <= my_rom(1567);
      when "011000100000" => q_unbuf <= my_rom(1568);
      when "011000100001" => q_unbuf <= my_rom(1569);
      when "011000100010" => q_unbuf <= my_rom(1570);
      when "011000100011" => q_unbuf <= my_rom(1571);
      when "011000100100" => q_unbuf <= my_rom(1572);
      when "011000100101" => q_unbuf <= my_rom(1573);
      when "011000100110" => q_unbuf <= my_rom(1574);
      when "011000100111" => q_unbuf <= my_rom(1575);
      when "011000101000" => q_unbuf <= my_rom(1576);
      when "011000101001" => q_unbuf <= my_rom(1577);
      when "011000101010" => q_unbuf <= my_rom(1578);
      when "011000101011" => q_unbuf <= my_rom(1579);
      when "011000101100" => q_unbuf <= my_rom(1580);
      when "011000101101" => q_unbuf <= my_rom(1581);
      when "011000101110" => q_unbuf <= my_rom(1582);
      when "011000101111" => q_unbuf <= my_rom(1583);
      when "011000110000" => q_unbuf <= my_rom(1584);
      when "011000110001" => q_unbuf <= my_rom(1585);
      when "011000110010" => q_unbuf <= my_rom(1586);
      when "011000110011" => q_unbuf <= my_rom(1587);
      when "011000110100" => q_unbuf <= my_rom(1588);
      when "011000110101" => q_unbuf <= my_rom(1589);
      when "011000110110" => q_unbuf <= my_rom(1590);
      when "011000110111" => q_unbuf <= my_rom(1591);
      when "011000111000" => q_unbuf <= my_rom(1592);
      when "011000111001" => q_unbuf <= my_rom(1593);
      when "011000111010" => q_unbuf <= my_rom(1594);
      when "011000111011" => q_unbuf <= my_rom(1595);
      when "011000111100" => q_unbuf <= my_rom(1596);
      when "011000111101" => q_unbuf <= my_rom(1597);
      when "011000111110" => q_unbuf <= my_rom(1598);
      when "011000111111" => q_unbuf <= my_rom(1599);
      when "011001000000" => q_unbuf <= my_rom(1600);
      when "011001000001" => q_unbuf <= my_rom(1601);
      when "011001000010" => q_unbuf <= my_rom(1602);
      when "011001000011" => q_unbuf <= my_rom(1603);
      when "011001000100" => q_unbuf <= my_rom(1604);
      when "011001000101" => q_unbuf <= my_rom(1605);
      when "011001000110" => q_unbuf <= my_rom(1606);
      when "011001000111" => q_unbuf <= my_rom(1607);
      when "011001001000" => q_unbuf <= my_rom(1608);
      when "011001001001" => q_unbuf <= my_rom(1609);
      when "011001001010" => q_unbuf <= my_rom(1610);
      when "011001001011" => q_unbuf <= my_rom(1611);
      when "011001001100" => q_unbuf <= my_rom(1612);
      when "011001001101" => q_unbuf <= my_rom(1613);
      when "011001001110" => q_unbuf <= my_rom(1614);
      when "011001001111" => q_unbuf <= my_rom(1615);
      when "011001010000" => q_unbuf <= my_rom(1616);
      when "011001010001" => q_unbuf <= my_rom(1617);
      when "011001010010" => q_unbuf <= my_rom(1618);
      when "011001010011" => q_unbuf <= my_rom(1619);
      when "011001010100" => q_unbuf <= my_rom(1620);
      when "011001010101" => q_unbuf <= my_rom(1621);
      when "011001010110" => q_unbuf <= my_rom(1622);
      when "011001010111" => q_unbuf <= my_rom(1623);
      when "011001011000" => q_unbuf <= my_rom(1624);
      when "011001011001" => q_unbuf <= my_rom(1625);
      when "011001011010" => q_unbuf <= my_rom(1626);
      when "011001011011" => q_unbuf <= my_rom(1627);
      when "011001011100" => q_unbuf <= my_rom(1628);
      when "011001011101" => q_unbuf <= my_rom(1629);
      when "011001011110" => q_unbuf <= my_rom(1630);
      when "011001011111" => q_unbuf <= my_rom(1631);
      when "011001100000" => q_unbuf <= my_rom(1632);
      when "011001100001" => q_unbuf <= my_rom(1633);
      when "011001100010" => q_unbuf <= my_rom(1634);
      when "011001100011" => q_unbuf <= my_rom(1635);
      when "011001100100" => q_unbuf <= my_rom(1636);
      when "011001100101" => q_unbuf <= my_rom(1637);
      when "011001100110" => q_unbuf <= my_rom(1638);
      when "011001100111" => q_unbuf <= my_rom(1639);
      when "011001101000" => q_unbuf <= my_rom(1640);
      when "011001101001" => q_unbuf <= my_rom(1641);
      when "011001101010" => q_unbuf <= my_rom(1642);
      when "011001101011" => q_unbuf <= my_rom(1643);
      when "011001101100" => q_unbuf <= my_rom(1644);
      when "011001101101" => q_unbuf <= my_rom(1645);
      when "011001101110" => q_unbuf <= my_rom(1646);
      when "011001101111" => q_unbuf <= my_rom(1647);
      when "011001110000" => q_unbuf <= my_rom(1648);
      when "011001110001" => q_unbuf <= my_rom(1649);
      when "011001110010" => q_unbuf <= my_rom(1650);
      when "011001110011" => q_unbuf <= my_rom(1651);
      when "011001110100" => q_unbuf <= my_rom(1652);
      when "011001110101" => q_unbuf <= my_rom(1653);
      when "011001110110" => q_unbuf <= my_rom(1654);
      when "011001110111" => q_unbuf <= my_rom(1655);
      when "011001111000" => q_unbuf <= my_rom(1656);
      when "011001111001" => q_unbuf <= my_rom(1657);
      when "011001111010" => q_unbuf <= my_rom(1658);
      when "011001111011" => q_unbuf <= my_rom(1659);
      when "011001111100" => q_unbuf <= my_rom(1660);
      when "011001111101" => q_unbuf <= my_rom(1661);
      when "011001111110" => q_unbuf <= my_rom(1662);
      when "011001111111" => q_unbuf <= my_rom(1663);
      when "011010000000" => q_unbuf <= my_rom(1664);
      when "011010000001" => q_unbuf <= my_rom(1665);
      when "011010000010" => q_unbuf <= my_rom(1666);
      when "011010000011" => q_unbuf <= my_rom(1667);
      when "011010000100" => q_unbuf <= my_rom(1668);
      when "011010000101" => q_unbuf <= my_rom(1669);
      when "011010000110" => q_unbuf <= my_rom(1670);
      when "011010000111" => q_unbuf <= my_rom(1671);
      when "011010001000" => q_unbuf <= my_rom(1672);
      when "011010001001" => q_unbuf <= my_rom(1673);
      when "011010001010" => q_unbuf <= my_rom(1674);
      when "011010001011" => q_unbuf <= my_rom(1675);
      when "011010001100" => q_unbuf <= my_rom(1676);
      when "011010001101" => q_unbuf <= my_rom(1677);
      when "011010001110" => q_unbuf <= my_rom(1678);
      when "011010001111" => q_unbuf <= my_rom(1679);
      when "011010010000" => q_unbuf <= my_rom(1680);
      when "011010010001" => q_unbuf <= my_rom(1681);
      when "011010010010" => q_unbuf <= my_rom(1682);
      when "011010010011" => q_unbuf <= my_rom(1683);
      when "011010010100" => q_unbuf <= my_rom(1684);
      when "011010010101" => q_unbuf <= my_rom(1685);
      when "011010010110" => q_unbuf <= my_rom(1686);
      when "011010010111" => q_unbuf <= my_rom(1687);
      when "011010011000" => q_unbuf <= my_rom(1688);
      when "011010011001" => q_unbuf <= my_rom(1689);
      when "011010011010" => q_unbuf <= my_rom(1690);
      when "011010011011" => q_unbuf <= my_rom(1691);
      when "011010011100" => q_unbuf <= my_rom(1692);
      when "011010011101" => q_unbuf <= my_rom(1693);
      when "011010011110" => q_unbuf <= my_rom(1694);
      when "011010011111" => q_unbuf <= my_rom(1695);
      when "011010100000" => q_unbuf <= my_rom(1696);
      when "011010100001" => q_unbuf <= my_rom(1697);
      when "011010100010" => q_unbuf <= my_rom(1698);
      when "011010100011" => q_unbuf <= my_rom(1699);
      when "011010100100" => q_unbuf <= my_rom(1700);
      when "011010100101" => q_unbuf <= my_rom(1701);
      when "011010100110" => q_unbuf <= my_rom(1702);
      when "011010100111" => q_unbuf <= my_rom(1703);
      when "011010101000" => q_unbuf <= my_rom(1704);
      when "011010101001" => q_unbuf <= my_rom(1705);
      when "011010101010" => q_unbuf <= my_rom(1706);
      when "011010101011" => q_unbuf <= my_rom(1707);
      when "011010101100" => q_unbuf <= my_rom(1708);
      when "011010101101" => q_unbuf <= my_rom(1709);
      when "011010101110" => q_unbuf <= my_rom(1710);
      when "011010101111" => q_unbuf <= my_rom(1711);
      when "011010110000" => q_unbuf <= my_rom(1712);
      when "011010110001" => q_unbuf <= my_rom(1713);
      when "011010110010" => q_unbuf <= my_rom(1714);
      when "011010110011" => q_unbuf <= my_rom(1715);
      when "011010110100" => q_unbuf <= my_rom(1716);
      when "011010110101" => q_unbuf <= my_rom(1717);
      when "011010110110" => q_unbuf <= my_rom(1718);
      when "011010110111" => q_unbuf <= my_rom(1719);
      when "011010111000" => q_unbuf <= my_rom(1720);
      when "011010111001" => q_unbuf <= my_rom(1721);
      when "011010111010" => q_unbuf <= my_rom(1722);
      when "011010111011" => q_unbuf <= my_rom(1723);
      when "011010111100" => q_unbuf <= my_rom(1724);
      when "011010111101" => q_unbuf <= my_rom(1725);
      when "011010111110" => q_unbuf <= my_rom(1726);
      when "011010111111" => q_unbuf <= my_rom(1727);
      when "011011000000" => q_unbuf <= my_rom(1728);
      when "011011000001" => q_unbuf <= my_rom(1729);
      when "011011000010" => q_unbuf <= my_rom(1730);
      when "011011000011" => q_unbuf <= my_rom(1731);
      when "011011000100" => q_unbuf <= my_rom(1732);
      when "011011000101" => q_unbuf <= my_rom(1733);
      when "011011000110" => q_unbuf <= my_rom(1734);
      when "011011000111" => q_unbuf <= my_rom(1735);
      when "011011001000" => q_unbuf <= my_rom(1736);
      when "011011001001" => q_unbuf <= my_rom(1737);
      when "011011001010" => q_unbuf <= my_rom(1738);
      when "011011001011" => q_unbuf <= my_rom(1739);
      when "011011001100" => q_unbuf <= my_rom(1740);
      when "011011001101" => q_unbuf <= my_rom(1741);
      when "011011001110" => q_unbuf <= my_rom(1742);
      when "011011001111" => q_unbuf <= my_rom(1743);
      when "011011010000" => q_unbuf <= my_rom(1744);
      when "011011010001" => q_unbuf <= my_rom(1745);
      when "011011010010" => q_unbuf <= my_rom(1746);
      when "011011010011" => q_unbuf <= my_rom(1747);
      when "011011010100" => q_unbuf <= my_rom(1748);
      when "011011010101" => q_unbuf <= my_rom(1749);
      when "011011010110" => q_unbuf <= my_rom(1750);
      when "011011010111" => q_unbuf <= my_rom(1751);
      when "011011011000" => q_unbuf <= my_rom(1752);
      when "011011011001" => q_unbuf <= my_rom(1753);
      when "011011011010" => q_unbuf <= my_rom(1754);
      when "011011011011" => q_unbuf <= my_rom(1755);
      when "011011011100" => q_unbuf <= my_rom(1756);
      when "011011011101" => q_unbuf <= my_rom(1757);
      when "011011011110" => q_unbuf <= my_rom(1758);
      when "011011011111" => q_unbuf <= my_rom(1759);
      when "011011100000" => q_unbuf <= my_rom(1760);
      when "011011100001" => q_unbuf <= my_rom(1761);
      when "011011100010" => q_unbuf <= my_rom(1762);
      when "011011100011" => q_unbuf <= my_rom(1763);
      when "011011100100" => q_unbuf <= my_rom(1764);
      when "011011100101" => q_unbuf <= my_rom(1765);
      when "011011100110" => q_unbuf <= my_rom(1766);
      when "011011100111" => q_unbuf <= my_rom(1767);
      when "011011101000" => q_unbuf <= my_rom(1768);
      when "011011101001" => q_unbuf <= my_rom(1769);
      when "011011101010" => q_unbuf <= my_rom(1770);
      when "011011101011" => q_unbuf <= my_rom(1771);
      when "011011101100" => q_unbuf <= my_rom(1772);
      when "011011101101" => q_unbuf <= my_rom(1773);
      when "011011101110" => q_unbuf <= my_rom(1774);
      when "011011101111" => q_unbuf <= my_rom(1775);
      when "011011110000" => q_unbuf <= my_rom(1776);
      when "011011110001" => q_unbuf <= my_rom(1777);
      when "011011110010" => q_unbuf <= my_rom(1778);
      when "011011110011" => q_unbuf <= my_rom(1779);
      when "011011110100" => q_unbuf <= my_rom(1780);
      when "011011110101" => q_unbuf <= my_rom(1781);
      when "011011110110" => q_unbuf <= my_rom(1782);
      when "011011110111" => q_unbuf <= my_rom(1783);
      when "011011111000" => q_unbuf <= my_rom(1784);
      when "011011111001" => q_unbuf <= my_rom(1785);
      when "011011111010" => q_unbuf <= my_rom(1786);
      when "011011111011" => q_unbuf <= my_rom(1787);
      when "011011111100" => q_unbuf <= my_rom(1788);
      when "011011111101" => q_unbuf <= my_rom(1789);
      when "011011111110" => q_unbuf <= my_rom(1790);
      when "011011111111" => q_unbuf <= my_rom(1791);
      when "011100000000" => q_unbuf <= my_rom(1792);
      when "011100000001" => q_unbuf <= my_rom(1793);
      when "011100000010" => q_unbuf <= my_rom(1794);
      when "011100000011" => q_unbuf <= my_rom(1795);
      when "011100000100" => q_unbuf <= my_rom(1796);
      when "011100000101" => q_unbuf <= my_rom(1797);
      when "011100000110" => q_unbuf <= my_rom(1798);
      when "011100000111" => q_unbuf <= my_rom(1799);
      when "011100001000" => q_unbuf <= my_rom(1800);
      when "011100001001" => q_unbuf <= my_rom(1801);
      when "011100001010" => q_unbuf <= my_rom(1802);
      when "011100001011" => q_unbuf <= my_rom(1803);
      when "011100001100" => q_unbuf <= my_rom(1804);
      when "011100001101" => q_unbuf <= my_rom(1805);
      when "011100001110" => q_unbuf <= my_rom(1806);
      when "011100001111" => q_unbuf <= my_rom(1807);
      when "011100010000" => q_unbuf <= my_rom(1808);
      when "011100010001" => q_unbuf <= my_rom(1809);
      when "011100010010" => q_unbuf <= my_rom(1810);
      when "011100010011" => q_unbuf <= my_rom(1811);
      when "011100010100" => q_unbuf <= my_rom(1812);
      when "011100010101" => q_unbuf <= my_rom(1813);
      when "011100010110" => q_unbuf <= my_rom(1814);
      when "011100010111" => q_unbuf <= my_rom(1815);
      when "011100011000" => q_unbuf <= my_rom(1816);
      when "011100011001" => q_unbuf <= my_rom(1817);
      when "011100011010" => q_unbuf <= my_rom(1818);
      when "011100011011" => q_unbuf <= my_rom(1819);
      when "011100011100" => q_unbuf <= my_rom(1820);
      when "011100011101" => q_unbuf <= my_rom(1821);
      when "011100011110" => q_unbuf <= my_rom(1822);
      when "011100011111" => q_unbuf <= my_rom(1823);
      when "011100100000" => q_unbuf <= my_rom(1824);
      when "011100100001" => q_unbuf <= my_rom(1825);
      when "011100100010" => q_unbuf <= my_rom(1826);
      when "011100100011" => q_unbuf <= my_rom(1827);
      when "011100100100" => q_unbuf <= my_rom(1828);
      when "011100100101" => q_unbuf <= my_rom(1829);
      when "011100100110" => q_unbuf <= my_rom(1830);
      when "011100100111" => q_unbuf <= my_rom(1831);
      when "011100101000" => q_unbuf <= my_rom(1832);
      when "011100101001" => q_unbuf <= my_rom(1833);
      when "011100101010" => q_unbuf <= my_rom(1834);
      when "011100101011" => q_unbuf <= my_rom(1835);
      when "011100101100" => q_unbuf <= my_rom(1836);
      when "011100101101" => q_unbuf <= my_rom(1837);
      when "011100101110" => q_unbuf <= my_rom(1838);
      when "011100101111" => q_unbuf <= my_rom(1839);
      when "011100110000" => q_unbuf <= my_rom(1840);
      when "011100110001" => q_unbuf <= my_rom(1841);
      when "011100110010" => q_unbuf <= my_rom(1842);
      when "011100110011" => q_unbuf <= my_rom(1843);
      when "011100110100" => q_unbuf <= my_rom(1844);
      when "011100110101" => q_unbuf <= my_rom(1845);
      when "011100110110" => q_unbuf <= my_rom(1846);
      when "011100110111" => q_unbuf <= my_rom(1847);
      when "011100111000" => q_unbuf <= my_rom(1848);
      when "011100111001" => q_unbuf <= my_rom(1849);
      when "011100111010" => q_unbuf <= my_rom(1850);
      when "011100111011" => q_unbuf <= my_rom(1851);
      when "011100111100" => q_unbuf <= my_rom(1852);
      when "011100111101" => q_unbuf <= my_rom(1853);
      when "011100111110" => q_unbuf <= my_rom(1854);
      when "011100111111" => q_unbuf <= my_rom(1855);
      when "011101000000" => q_unbuf <= my_rom(1856);
      when "011101000001" => q_unbuf <= my_rom(1857);
      when "011101000010" => q_unbuf <= my_rom(1858);
      when "011101000011" => q_unbuf <= my_rom(1859);
      when "011101000100" => q_unbuf <= my_rom(1860);
      when "011101000101" => q_unbuf <= my_rom(1861);
      when "011101000110" => q_unbuf <= my_rom(1862);
      when "011101000111" => q_unbuf <= my_rom(1863);
      when "011101001000" => q_unbuf <= my_rom(1864);
      when "011101001001" => q_unbuf <= my_rom(1865);
      when "011101001010" => q_unbuf <= my_rom(1866);
      when "011101001011" => q_unbuf <= my_rom(1867);
      when "011101001100" => q_unbuf <= my_rom(1868);
      when "011101001101" => q_unbuf <= my_rom(1869);
      when "011101001110" => q_unbuf <= my_rom(1870);
      when "011101001111" => q_unbuf <= my_rom(1871);
      when "011101010000" => q_unbuf <= my_rom(1872);
      when "011101010001" => q_unbuf <= my_rom(1873);
      when "011101010010" => q_unbuf <= my_rom(1874);
      when "011101010011" => q_unbuf <= my_rom(1875);
      when "011101010100" => q_unbuf <= my_rom(1876);
      when "011101010101" => q_unbuf <= my_rom(1877);
      when "011101010110" => q_unbuf <= my_rom(1878);
      when "011101010111" => q_unbuf <= my_rom(1879);
      when "011101011000" => q_unbuf <= my_rom(1880);
      when "011101011001" => q_unbuf <= my_rom(1881);
      when "011101011010" => q_unbuf <= my_rom(1882);
      when "011101011011" => q_unbuf <= my_rom(1883);
      when "011101011100" => q_unbuf <= my_rom(1884);
      when "011101011101" => q_unbuf <= my_rom(1885);
      when "011101011110" => q_unbuf <= my_rom(1886);
      when "011101011111" => q_unbuf <= my_rom(1887);
      when "011101100000" => q_unbuf <= my_rom(1888);
      when "011101100001" => q_unbuf <= my_rom(1889);
      when "011101100010" => q_unbuf <= my_rom(1890);
      when "011101100011" => q_unbuf <= my_rom(1891);
      when "011101100100" => q_unbuf <= my_rom(1892);
      when "011101100101" => q_unbuf <= my_rom(1893);
      when "011101100110" => q_unbuf <= my_rom(1894);
      when "011101100111" => q_unbuf <= my_rom(1895);
      when "011101101000" => q_unbuf <= my_rom(1896);
      when "011101101001" => q_unbuf <= my_rom(1897);
      when "011101101010" => q_unbuf <= my_rom(1898);
      when "011101101011" => q_unbuf <= my_rom(1899);
      when "011101101100" => q_unbuf <= my_rom(1900);
      when "011101101101" => q_unbuf <= my_rom(1901);
      when "011101101110" => q_unbuf <= my_rom(1902);
      when "011101101111" => q_unbuf <= my_rom(1903);
      when "011101110000" => q_unbuf <= my_rom(1904);
      when "011101110001" => q_unbuf <= my_rom(1905);
      when "011101110010" => q_unbuf <= my_rom(1906);
      when "011101110011" => q_unbuf <= my_rom(1907);
      when "011101110100" => q_unbuf <= my_rom(1908);
      when "011101110101" => q_unbuf <= my_rom(1909);
      when "011101110110" => q_unbuf <= my_rom(1910);
      when "011101110111" => q_unbuf <= my_rom(1911);
      when "011101111000" => q_unbuf <= my_rom(1912);
      when "011101111001" => q_unbuf <= my_rom(1913);
      when "011101111010" => q_unbuf <= my_rom(1914);
      when "011101111011" => q_unbuf <= my_rom(1915);
      when "011101111100" => q_unbuf <= my_rom(1916);
      when "011101111101" => q_unbuf <= my_rom(1917);
      when "011101111110" => q_unbuf <= my_rom(1918);
      when "011101111111" => q_unbuf <= my_rom(1919);
      when "011110000000" => q_unbuf <= my_rom(1920);
      when "011110000001" => q_unbuf <= my_rom(1921);
      when "011110000010" => q_unbuf <= my_rom(1922);
      when "011110000011" => q_unbuf <= my_rom(1923);
      when "011110000100" => q_unbuf <= my_rom(1924);
      when "011110000101" => q_unbuf <= my_rom(1925);
      when "011110000110" => q_unbuf <= my_rom(1926);
      when "011110000111" => q_unbuf <= my_rom(1927);
      when "011110001000" => q_unbuf <= my_rom(1928);
      when "011110001001" => q_unbuf <= my_rom(1929);
      when "011110001010" => q_unbuf <= my_rom(1930);
      when "011110001011" => q_unbuf <= my_rom(1931);
      when "011110001100" => q_unbuf <= my_rom(1932);
      when "011110001101" => q_unbuf <= my_rom(1933);
      when "011110001110" => q_unbuf <= my_rom(1934);
      when "011110001111" => q_unbuf <= my_rom(1935);
      when "011110010000" => q_unbuf <= my_rom(1936);
      when "011110010001" => q_unbuf <= my_rom(1937);
      when "011110010010" => q_unbuf <= my_rom(1938);
      when "011110010011" => q_unbuf <= my_rom(1939);
      when "011110010100" => q_unbuf <= my_rom(1940);
      when "011110010101" => q_unbuf <= my_rom(1941);
      when "011110010110" => q_unbuf <= my_rom(1942);
      when "011110010111" => q_unbuf <= my_rom(1943);
      when "011110011000" => q_unbuf <= my_rom(1944);
      when "011110011001" => q_unbuf <= my_rom(1945);
      when "011110011010" => q_unbuf <= my_rom(1946);
      when "011110011011" => q_unbuf <= my_rom(1947);
      when "011110011100" => q_unbuf <= my_rom(1948);
      when "011110011101" => q_unbuf <= my_rom(1949);
      when "011110011110" => q_unbuf <= my_rom(1950);
      when "011110011111" => q_unbuf <= my_rom(1951);
      when "011110100000" => q_unbuf <= my_rom(1952);
      when "011110100001" => q_unbuf <= my_rom(1953);
      when "011110100010" => q_unbuf <= my_rom(1954);
      when "011110100011" => q_unbuf <= my_rom(1955);
      when "011110100100" => q_unbuf <= my_rom(1956);
      when "011110100101" => q_unbuf <= my_rom(1957);
      when "011110100110" => q_unbuf <= my_rom(1958);
      when "011110100111" => q_unbuf <= my_rom(1959);
      when "011110101000" => q_unbuf <= my_rom(1960);
      when "011110101001" => q_unbuf <= my_rom(1961);
      when "011110101010" => q_unbuf <= my_rom(1962);
      when "011110101011" => q_unbuf <= my_rom(1963);
      when "011110101100" => q_unbuf <= my_rom(1964);
      when "011110101101" => q_unbuf <= my_rom(1965);
      when "011110101110" => q_unbuf <= my_rom(1966);
      when "011110101111" => q_unbuf <= my_rom(1967);
      when "011110110000" => q_unbuf <= my_rom(1968);
      when "011110110001" => q_unbuf <= my_rom(1969);
      when "011110110010" => q_unbuf <= my_rom(1970);
      when "011110110011" => q_unbuf <= my_rom(1971);
      when "011110110100" => q_unbuf <= my_rom(1972);
      when "011110110101" => q_unbuf <= my_rom(1973);
      when "011110110110" => q_unbuf <= my_rom(1974);
      when "011110110111" => q_unbuf <= my_rom(1975);
      when "011110111000" => q_unbuf <= my_rom(1976);
      when "011110111001" => q_unbuf <= my_rom(1977);
      when "011110111010" => q_unbuf <= my_rom(1978);
      when "011110111011" => q_unbuf <= my_rom(1979);
      when "011110111100" => q_unbuf <= my_rom(1980);
      when "011110111101" => q_unbuf <= my_rom(1981);
      when "011110111110" => q_unbuf <= my_rom(1982);
      when "011110111111" => q_unbuf <= my_rom(1983);
      when "011111000000" => q_unbuf <= my_rom(1984);
      when "011111000001" => q_unbuf <= my_rom(1985);
      when "011111000010" => q_unbuf <= my_rom(1986);
      when "011111000011" => q_unbuf <= my_rom(1987);
      when "011111000100" => q_unbuf <= my_rom(1988);
      when "011111000101" => q_unbuf <= my_rom(1989);
      when "011111000110" => q_unbuf <= my_rom(1990);
      when "011111000111" => q_unbuf <= my_rom(1991);
      when "011111001000" => q_unbuf <= my_rom(1992);
      when "011111001001" => q_unbuf <= my_rom(1993);
      when "011111001010" => q_unbuf <= my_rom(1994);
      when "011111001011" => q_unbuf <= my_rom(1995);
      when "011111001100" => q_unbuf <= my_rom(1996);
      when "011111001101" => q_unbuf <= my_rom(1997);
      when "011111001110" => q_unbuf <= my_rom(1998);
      when "011111001111" => q_unbuf <= my_rom(1999);
      when "011111010000" => q_unbuf <= my_rom(2000);
      when "011111010001" => q_unbuf <= my_rom(2001);
      when "011111010010" => q_unbuf <= my_rom(2002);
      when "011111010011" => q_unbuf <= my_rom(2003);
      when "011111010100" => q_unbuf <= my_rom(2004);
      when "011111010101" => q_unbuf <= my_rom(2005);
      when "011111010110" => q_unbuf <= my_rom(2006);
      when "011111010111" => q_unbuf <= my_rom(2007);
      when "011111011000" => q_unbuf <= my_rom(2008);
      when "011111011001" => q_unbuf <= my_rom(2009);
      when "011111011010" => q_unbuf <= my_rom(2010);
      when "011111011011" => q_unbuf <= my_rom(2011);
      when "011111011100" => q_unbuf <= my_rom(2012);
      when "011111011101" => q_unbuf <= my_rom(2013);
      when "011111011110" => q_unbuf <= my_rom(2014);
      when "011111011111" => q_unbuf <= my_rom(2015);
      when "011111100000" => q_unbuf <= my_rom(2016);
      when "011111100001" => q_unbuf <= my_rom(2017);
      when "011111100010" => q_unbuf <= my_rom(2018);
      when "011111100011" => q_unbuf <= my_rom(2019);
      when "011111100100" => q_unbuf <= my_rom(2020);
      when "011111100101" => q_unbuf <= my_rom(2021);
      when "011111100110" => q_unbuf <= my_rom(2022);
      when "011111100111" => q_unbuf <= my_rom(2023);
      when "011111101000" => q_unbuf <= my_rom(2024);
      when "011111101001" => q_unbuf <= my_rom(2025);
      when "011111101010" => q_unbuf <= my_rom(2026);
      when "011111101011" => q_unbuf <= my_rom(2027);
      when "011111101100" => q_unbuf <= my_rom(2028);
      when "011111101101" => q_unbuf <= my_rom(2029);
      when "011111101110" => q_unbuf <= my_rom(2030);
      when "011111101111" => q_unbuf <= my_rom(2031);
      when "011111110000" => q_unbuf <= my_rom(2032);
      when "011111110001" => q_unbuf <= my_rom(2033);
      when "011111110010" => q_unbuf <= my_rom(2034);
      when "011111110011" => q_unbuf <= my_rom(2035);
      when "011111110100" => q_unbuf <= my_rom(2036);
      when "011111110101" => q_unbuf <= my_rom(2037);
      when "011111110110" => q_unbuf <= my_rom(2038);
      when "011111110111" => q_unbuf <= my_rom(2039);
      when "011111111000" => q_unbuf <= my_rom(2040);
      when "011111111001" => q_unbuf <= my_rom(2041);
      when "011111111010" => q_unbuf <= my_rom(2042);
      when "011111111011" => q_unbuf <= my_rom(2043);
      when "011111111100" => q_unbuf <= my_rom(2044);
      when "011111111101" => q_unbuf <= my_rom(2045);
      when "011111111110" => q_unbuf <= my_rom(2046);
      when "011111111111" => q_unbuf <= my_rom(2047);
      when "100000000000" => q_unbuf <= my_rom(2048);
      when "100000000001" => q_unbuf <= my_rom(2049);
      when "100000000010" => q_unbuf <= my_rom(2050);
      when "100000000011" => q_unbuf <= my_rom(2051);
      when "100000000100" => q_unbuf <= my_rom(2052);
      when "100000000101" => q_unbuf <= my_rom(2053);
      when "100000000110" => q_unbuf <= my_rom(2054);
      when "100000000111" => q_unbuf <= my_rom(2055);
      when "100000001000" => q_unbuf <= my_rom(2056);
      when "100000001001" => q_unbuf <= my_rom(2057);
      when "100000001010" => q_unbuf <= my_rom(2058);
      when "100000001011" => q_unbuf <= my_rom(2059);
      when "100000001100" => q_unbuf <= my_rom(2060);
      when "100000001101" => q_unbuf <= my_rom(2061);
      when "100000001110" => q_unbuf <= my_rom(2062);
      when "100000001111" => q_unbuf <= my_rom(2063);
      when "100000010000" => q_unbuf <= my_rom(2064);
      when "100000010001" => q_unbuf <= my_rom(2065);
      when "100000010010" => q_unbuf <= my_rom(2066);
      when "100000010011" => q_unbuf <= my_rom(2067);
      when "100000010100" => q_unbuf <= my_rom(2068);
      when "100000010101" => q_unbuf <= my_rom(2069);
      when "100000010110" => q_unbuf <= my_rom(2070);
      when "100000010111" => q_unbuf <= my_rom(2071);
      when "100000011000" => q_unbuf <= my_rom(2072);
      when "100000011001" => q_unbuf <= my_rom(2073);
      when "100000011010" => q_unbuf <= my_rom(2074);
      when "100000011011" => q_unbuf <= my_rom(2075);
      when "100000011100" => q_unbuf <= my_rom(2076);
      when "100000011101" => q_unbuf <= my_rom(2077);
      when "100000011110" => q_unbuf <= my_rom(2078);
      when "100000011111" => q_unbuf <= my_rom(2079);
      when "100000100000" => q_unbuf <= my_rom(2080);
      when "100000100001" => q_unbuf <= my_rom(2081);
      when "100000100010" => q_unbuf <= my_rom(2082);
      when "100000100011" => q_unbuf <= my_rom(2083);
      when "100000100100" => q_unbuf <= my_rom(2084);
      when "100000100101" => q_unbuf <= my_rom(2085);
      when "100000100110" => q_unbuf <= my_rom(2086);
      when "100000100111" => q_unbuf <= my_rom(2087);
      when "100000101000" => q_unbuf <= my_rom(2088);
      when "100000101001" => q_unbuf <= my_rom(2089);
      when "100000101010" => q_unbuf <= my_rom(2090);
      when "100000101011" => q_unbuf <= my_rom(2091);
      when "100000101100" => q_unbuf <= my_rom(2092);
      when "100000101101" => q_unbuf <= my_rom(2093);
      when "100000101110" => q_unbuf <= my_rom(2094);
      when "100000101111" => q_unbuf <= my_rom(2095);
      when "100000110000" => q_unbuf <= my_rom(2096);
      when "100000110001" => q_unbuf <= my_rom(2097);
      when "100000110010" => q_unbuf <= my_rom(2098);
      when "100000110011" => q_unbuf <= my_rom(2099);
      when "100000110100" => q_unbuf <= my_rom(2100);
      when "100000110101" => q_unbuf <= my_rom(2101);
      when "100000110110" => q_unbuf <= my_rom(2102);
      when "100000110111" => q_unbuf <= my_rom(2103);
      when "100000111000" => q_unbuf <= my_rom(2104);
      when "100000111001" => q_unbuf <= my_rom(2105);
      when "100000111010" => q_unbuf <= my_rom(2106);
      when "100000111011" => q_unbuf <= my_rom(2107);
      when "100000111100" => q_unbuf <= my_rom(2108);
      when "100000111101" => q_unbuf <= my_rom(2109);
      when "100000111110" => q_unbuf <= my_rom(2110);
      when "100000111111" => q_unbuf <= my_rom(2111);
      when "100001000000" => q_unbuf <= my_rom(2112);
      when "100001000001" => q_unbuf <= my_rom(2113);
      when "100001000010" => q_unbuf <= my_rom(2114);
      when "100001000011" => q_unbuf <= my_rom(2115);
      when "100001000100" => q_unbuf <= my_rom(2116);
      when "100001000101" => q_unbuf <= my_rom(2117);
      when "100001000110" => q_unbuf <= my_rom(2118);
      when "100001000111" => q_unbuf <= my_rom(2119);
      when "100001001000" => q_unbuf <= my_rom(2120);
      when "100001001001" => q_unbuf <= my_rom(2121);
      when "100001001010" => q_unbuf <= my_rom(2122);
      when "100001001011" => q_unbuf <= my_rom(2123);
      when "100001001100" => q_unbuf <= my_rom(2124);
      when "100001001101" => q_unbuf <= my_rom(2125);
      when "100001001110" => q_unbuf <= my_rom(2126);
      when "100001001111" => q_unbuf <= my_rom(2127);
      when "100001010000" => q_unbuf <= my_rom(2128);
      when "100001010001" => q_unbuf <= my_rom(2129);
      when "100001010010" => q_unbuf <= my_rom(2130);
      when "100001010011" => q_unbuf <= my_rom(2131);
      when "100001010100" => q_unbuf <= my_rom(2132);
      when "100001010101" => q_unbuf <= my_rom(2133);
      when "100001010110" => q_unbuf <= my_rom(2134);
      when "100001010111" => q_unbuf <= my_rom(2135);
      when "100001011000" => q_unbuf <= my_rom(2136);
      when "100001011001" => q_unbuf <= my_rom(2137);
      when "100001011010" => q_unbuf <= my_rom(2138);
      when "100001011011" => q_unbuf <= my_rom(2139);
      when "100001011100" => q_unbuf <= my_rom(2140);
      when "100001011101" => q_unbuf <= my_rom(2141);
      when "100001011110" => q_unbuf <= my_rom(2142);
      when "100001011111" => q_unbuf <= my_rom(2143);
      when "100001100000" => q_unbuf <= my_rom(2144);
      when "100001100001" => q_unbuf <= my_rom(2145);
      when "100001100010" => q_unbuf <= my_rom(2146);
      when "100001100011" => q_unbuf <= my_rom(2147);
      when "100001100100" => q_unbuf <= my_rom(2148);
      when "100001100101" => q_unbuf <= my_rom(2149);
      when "100001100110" => q_unbuf <= my_rom(2150);
      when "100001100111" => q_unbuf <= my_rom(2151);
      when "100001101000" => q_unbuf <= my_rom(2152);
      when "100001101001" => q_unbuf <= my_rom(2153);
      when "100001101010" => q_unbuf <= my_rom(2154);
      when "100001101011" => q_unbuf <= my_rom(2155);
      when "100001101100" => q_unbuf <= my_rom(2156);
      when "100001101101" => q_unbuf <= my_rom(2157);
      when "100001101110" => q_unbuf <= my_rom(2158);
      when "100001101111" => q_unbuf <= my_rom(2159);
      when "100001110000" => q_unbuf <= my_rom(2160);
      when "100001110001" => q_unbuf <= my_rom(2161);
      when "100001110010" => q_unbuf <= my_rom(2162);
      when "100001110011" => q_unbuf <= my_rom(2163);
      when "100001110100" => q_unbuf <= my_rom(2164);
      when "100001110101" => q_unbuf <= my_rom(2165);
      when "100001110110" => q_unbuf <= my_rom(2166);
      when "100001110111" => q_unbuf <= my_rom(2167);
      when "100001111000" => q_unbuf <= my_rom(2168);
      when "100001111001" => q_unbuf <= my_rom(2169);
      when "100001111010" => q_unbuf <= my_rom(2170);
      when "100001111011" => q_unbuf <= my_rom(2171);
      when "100001111100" => q_unbuf <= my_rom(2172);
      when "100001111101" => q_unbuf <= my_rom(2173);
      when "100001111110" => q_unbuf <= my_rom(2174);
      when "100001111111" => q_unbuf <= my_rom(2175);
      when "100010000000" => q_unbuf <= my_rom(2176);
      when "100010000001" => q_unbuf <= my_rom(2177);
      when "100010000010" => q_unbuf <= my_rom(2178);
      when "100010000011" => q_unbuf <= my_rom(2179);
      when "100010000100" => q_unbuf <= my_rom(2180);
      when "100010000101" => q_unbuf <= my_rom(2181);
      when "100010000110" => q_unbuf <= my_rom(2182);
      when "100010000111" => q_unbuf <= my_rom(2183);
      when "100010001000" => q_unbuf <= my_rom(2184);
      when "100010001001" => q_unbuf <= my_rom(2185);
      when "100010001010" => q_unbuf <= my_rom(2186);
      when "100010001011" => q_unbuf <= my_rom(2187);
      when "100010001100" => q_unbuf <= my_rom(2188);
      when "100010001101" => q_unbuf <= my_rom(2189);
      when "100010001110" => q_unbuf <= my_rom(2190);
      when "100010001111" => q_unbuf <= my_rom(2191);
      when "100010010000" => q_unbuf <= my_rom(2192);
      when "100010010001" => q_unbuf <= my_rom(2193);
      when "100010010010" => q_unbuf <= my_rom(2194);
      when "100010010011" => q_unbuf <= my_rom(2195);
      when "100010010100" => q_unbuf <= my_rom(2196);
      when "100010010101" => q_unbuf <= my_rom(2197);
      when "100010010110" => q_unbuf <= my_rom(2198);
      when "100010010111" => q_unbuf <= my_rom(2199);
      when "100010011000" => q_unbuf <= my_rom(2200);
      when "100010011001" => q_unbuf <= my_rom(2201);
      when "100010011010" => q_unbuf <= my_rom(2202);
      when "100010011011" => q_unbuf <= my_rom(2203);
      when "100010011100" => q_unbuf <= my_rom(2204);
      when "100010011101" => q_unbuf <= my_rom(2205);
      when "100010011110" => q_unbuf <= my_rom(2206);
      when "100010011111" => q_unbuf <= my_rom(2207);
      when "100010100000" => q_unbuf <= my_rom(2208);
      when "100010100001" => q_unbuf <= my_rom(2209);
      when "100010100010" => q_unbuf <= my_rom(2210);
      when "100010100011" => q_unbuf <= my_rom(2211);
      when "100010100100" => q_unbuf <= my_rom(2212);
      when "100010100101" => q_unbuf <= my_rom(2213);
      when "100010100110" => q_unbuf <= my_rom(2214);
      when "100010100111" => q_unbuf <= my_rom(2215);
      when "100010101000" => q_unbuf <= my_rom(2216);
      when "100010101001" => q_unbuf <= my_rom(2217);
      when "100010101010" => q_unbuf <= my_rom(2218);
      when "100010101011" => q_unbuf <= my_rom(2219);
      when "100010101100" => q_unbuf <= my_rom(2220);
      when "100010101101" => q_unbuf <= my_rom(2221);
      when "100010101110" => q_unbuf <= my_rom(2222);
      when "100010101111" => q_unbuf <= my_rom(2223);
      when "100010110000" => q_unbuf <= my_rom(2224);
      when "100010110001" => q_unbuf <= my_rom(2225);
      when "100010110010" => q_unbuf <= my_rom(2226);
      when "100010110011" => q_unbuf <= my_rom(2227);
      when "100010110100" => q_unbuf <= my_rom(2228);
      when "100010110101" => q_unbuf <= my_rom(2229);
      when "100010110110" => q_unbuf <= my_rom(2230);
      when "100010110111" => q_unbuf <= my_rom(2231);
      when "100010111000" => q_unbuf <= my_rom(2232);
      when "100010111001" => q_unbuf <= my_rom(2233);
      when "100010111010" => q_unbuf <= my_rom(2234);
      when "100010111011" => q_unbuf <= my_rom(2235);
      when "100010111100" => q_unbuf <= my_rom(2236);
      when "100010111101" => q_unbuf <= my_rom(2237);
      when "100010111110" => q_unbuf <= my_rom(2238);
      when "100010111111" => q_unbuf <= my_rom(2239);
      when "100011000000" => q_unbuf <= my_rom(2240);
      when "100011000001" => q_unbuf <= my_rom(2241);
      when "100011000010" => q_unbuf <= my_rom(2242);
      when "100011000011" => q_unbuf <= my_rom(2243);
      when "100011000100" => q_unbuf <= my_rom(2244);
      when "100011000101" => q_unbuf <= my_rom(2245);
      when "100011000110" => q_unbuf <= my_rom(2246);
      when "100011000111" => q_unbuf <= my_rom(2247);
      when "100011001000" => q_unbuf <= my_rom(2248);
      when "100011001001" => q_unbuf <= my_rom(2249);
      when "100011001010" => q_unbuf <= my_rom(2250);
      when "100011001011" => q_unbuf <= my_rom(2251);
      when "100011001100" => q_unbuf <= my_rom(2252);
      when "100011001101" => q_unbuf <= my_rom(2253);
      when "100011001110" => q_unbuf <= my_rom(2254);
      when "100011001111" => q_unbuf <= my_rom(2255);
      when "100011010000" => q_unbuf <= my_rom(2256);
      when "100011010001" => q_unbuf <= my_rom(2257);
      when "100011010010" => q_unbuf <= my_rom(2258);
      when "100011010011" => q_unbuf <= my_rom(2259);
      when "100011010100" => q_unbuf <= my_rom(2260);
      when "100011010101" => q_unbuf <= my_rom(2261);
      when "100011010110" => q_unbuf <= my_rom(2262);
      when "100011010111" => q_unbuf <= my_rom(2263);
      when "100011011000" => q_unbuf <= my_rom(2264);
      when "100011011001" => q_unbuf <= my_rom(2265);
      when "100011011010" => q_unbuf <= my_rom(2266);
      when "100011011011" => q_unbuf <= my_rom(2267);
      when "100011011100" => q_unbuf <= my_rom(2268);
      when "100011011101" => q_unbuf <= my_rom(2269);
      when "100011011110" => q_unbuf <= my_rom(2270);
      when "100011011111" => q_unbuf <= my_rom(2271);
      when "100011100000" => q_unbuf <= my_rom(2272);
      when "100011100001" => q_unbuf <= my_rom(2273);
      when "100011100010" => q_unbuf <= my_rom(2274);
      when "100011100011" => q_unbuf <= my_rom(2275);
      when "100011100100" => q_unbuf <= my_rom(2276);
      when "100011100101" => q_unbuf <= my_rom(2277);
      when "100011100110" => q_unbuf <= my_rom(2278);
      when "100011100111" => q_unbuf <= my_rom(2279);
      when "100011101000" => q_unbuf <= my_rom(2280);
      when "100011101001" => q_unbuf <= my_rom(2281);
      when "100011101010" => q_unbuf <= my_rom(2282);
      when "100011101011" => q_unbuf <= my_rom(2283);
      when "100011101100" => q_unbuf <= my_rom(2284);
      when "100011101101" => q_unbuf <= my_rom(2285);
      when "100011101110" => q_unbuf <= my_rom(2286);
      when "100011101111" => q_unbuf <= my_rom(2287);
      when "100011110000" => q_unbuf <= my_rom(2288);
      when "100011110001" => q_unbuf <= my_rom(2289);
      when "100011110010" => q_unbuf <= my_rom(2290);
      when "100011110011" => q_unbuf <= my_rom(2291);
      when "100011110100" => q_unbuf <= my_rom(2292);
      when "100011110101" => q_unbuf <= my_rom(2293);
      when "100011110110" => q_unbuf <= my_rom(2294);
      when "100011110111" => q_unbuf <= my_rom(2295);
      when "100011111000" => q_unbuf <= my_rom(2296);
      when "100011111001" => q_unbuf <= my_rom(2297);
      when "100011111010" => q_unbuf <= my_rom(2298);
      when "100011111011" => q_unbuf <= my_rom(2299);
      when "100011111100" => q_unbuf <= my_rom(2300);
      when "100011111101" => q_unbuf <= my_rom(2301);
      when "100011111110" => q_unbuf <= my_rom(2302);
      when "100011111111" => q_unbuf <= my_rom(2303);
      when "100100000000" => q_unbuf <= my_rom(2304);
      when "100100000001" => q_unbuf <= my_rom(2305);
      when "100100000010" => q_unbuf <= my_rom(2306);
      when "100100000011" => q_unbuf <= my_rom(2307);
      when "100100000100" => q_unbuf <= my_rom(2308);
      when "100100000101" => q_unbuf <= my_rom(2309);
      when "100100000110" => q_unbuf <= my_rom(2310);
      when "100100000111" => q_unbuf <= my_rom(2311);
      when "100100001000" => q_unbuf <= my_rom(2312);
      when "100100001001" => q_unbuf <= my_rom(2313);
      when "100100001010" => q_unbuf <= my_rom(2314);
      when "100100001011" => q_unbuf <= my_rom(2315);
      when "100100001100" => q_unbuf <= my_rom(2316);
      when "100100001101" => q_unbuf <= my_rom(2317);
      when "100100001110" => q_unbuf <= my_rom(2318);
      when "100100001111" => q_unbuf <= my_rom(2319);
      when "100100010000" => q_unbuf <= my_rom(2320);
      when "100100010001" => q_unbuf <= my_rom(2321);
      when "100100010010" => q_unbuf <= my_rom(2322);
      when "100100010011" => q_unbuf <= my_rom(2323);
      when "100100010100" => q_unbuf <= my_rom(2324);
      when "100100010101" => q_unbuf <= my_rom(2325);
      when "100100010110" => q_unbuf <= my_rom(2326);
      when "100100010111" => q_unbuf <= my_rom(2327);
      when "100100011000" => q_unbuf <= my_rom(2328);
      when "100100011001" => q_unbuf <= my_rom(2329);
      when "100100011010" => q_unbuf <= my_rom(2330);
      when "100100011011" => q_unbuf <= my_rom(2331);
      when "100100011100" => q_unbuf <= my_rom(2332);
      when "100100011101" => q_unbuf <= my_rom(2333);
      when "100100011110" => q_unbuf <= my_rom(2334);
      when "100100011111" => q_unbuf <= my_rom(2335);
      when "100100100000" => q_unbuf <= my_rom(2336);
      when "100100100001" => q_unbuf <= my_rom(2337);
      when "100100100010" => q_unbuf <= my_rom(2338);
      when "100100100011" => q_unbuf <= my_rom(2339);
      when "100100100100" => q_unbuf <= my_rom(2340);
      when "100100100101" => q_unbuf <= my_rom(2341);
      when "100100100110" => q_unbuf <= my_rom(2342);
      when "100100100111" => q_unbuf <= my_rom(2343);
      when "100100101000" => q_unbuf <= my_rom(2344);
      when "100100101001" => q_unbuf <= my_rom(2345);
      when "100100101010" => q_unbuf <= my_rom(2346);
      when "100100101011" => q_unbuf <= my_rom(2347);
      when "100100101100" => q_unbuf <= my_rom(2348);
      when "100100101101" => q_unbuf <= my_rom(2349);
      when "100100101110" => q_unbuf <= my_rom(2350);
      when "100100101111" => q_unbuf <= my_rom(2351);
      when "100100110000" => q_unbuf <= my_rom(2352);
      when "100100110001" => q_unbuf <= my_rom(2353);
      when "100100110010" => q_unbuf <= my_rom(2354);
      when "100100110011" => q_unbuf <= my_rom(2355);
      when "100100110100" => q_unbuf <= my_rom(2356);
      when "100100110101" => q_unbuf <= my_rom(2357);
      when "100100110110" => q_unbuf <= my_rom(2358);
      when "100100110111" => q_unbuf <= my_rom(2359);
      when "100100111000" => q_unbuf <= my_rom(2360);
      when "100100111001" => q_unbuf <= my_rom(2361);
      when "100100111010" => q_unbuf <= my_rom(2362);
      when "100100111011" => q_unbuf <= my_rom(2363);
      when "100100111100" => q_unbuf <= my_rom(2364);
      when "100100111101" => q_unbuf <= my_rom(2365);
      when "100100111110" => q_unbuf <= my_rom(2366);
      when "100100111111" => q_unbuf <= my_rom(2367);
      when "100101000000" => q_unbuf <= my_rom(2368);
      when "100101000001" => q_unbuf <= my_rom(2369);
      when "100101000010" => q_unbuf <= my_rom(2370);
      when "100101000011" => q_unbuf <= my_rom(2371);
      when "100101000100" => q_unbuf <= my_rom(2372);
      when "100101000101" => q_unbuf <= my_rom(2373);
      when "100101000110" => q_unbuf <= my_rom(2374);
      when "100101000111" => q_unbuf <= my_rom(2375);
      when "100101001000" => q_unbuf <= my_rom(2376);
      when "100101001001" => q_unbuf <= my_rom(2377);
      when "100101001010" => q_unbuf <= my_rom(2378);
      when "100101001011" => q_unbuf <= my_rom(2379);
      when "100101001100" => q_unbuf <= my_rom(2380);
      when "100101001101" => q_unbuf <= my_rom(2381);
      when "100101001110" => q_unbuf <= my_rom(2382);
      when "100101001111" => q_unbuf <= my_rom(2383);
      when "100101010000" => q_unbuf <= my_rom(2384);
      when "100101010001" => q_unbuf <= my_rom(2385);
      when "100101010010" => q_unbuf <= my_rom(2386);
      when "100101010011" => q_unbuf <= my_rom(2387);
      when "100101010100" => q_unbuf <= my_rom(2388);
      when "100101010101" => q_unbuf <= my_rom(2389);
      when "100101010110" => q_unbuf <= my_rom(2390);
      when "100101010111" => q_unbuf <= my_rom(2391);
      when "100101011000" => q_unbuf <= my_rom(2392);
      when "100101011001" => q_unbuf <= my_rom(2393);
      when "100101011010" => q_unbuf <= my_rom(2394);
      when "100101011011" => q_unbuf <= my_rom(2395);
      when "100101011100" => q_unbuf <= my_rom(2396);
      when "100101011101" => q_unbuf <= my_rom(2397);
      when "100101011110" => q_unbuf <= my_rom(2398);
      when "100101011111" => q_unbuf <= my_rom(2399);
      when "100101100000" => q_unbuf <= my_rom(2400);
      when "100101100001" => q_unbuf <= my_rom(2401);
      when "100101100010" => q_unbuf <= my_rom(2402);
      when "100101100011" => q_unbuf <= my_rom(2403);
      when "100101100100" => q_unbuf <= my_rom(2404);
      when "100101100101" => q_unbuf <= my_rom(2405);
      when "100101100110" => q_unbuf <= my_rom(2406);
      when "100101100111" => q_unbuf <= my_rom(2407);
      when "100101101000" => q_unbuf <= my_rom(2408);
      when "100101101001" => q_unbuf <= my_rom(2409);
      when "100101101010" => q_unbuf <= my_rom(2410);
      when "100101101011" => q_unbuf <= my_rom(2411);
      when "100101101100" => q_unbuf <= my_rom(2412);
      when "100101101101" => q_unbuf <= my_rom(2413);
      when "100101101110" => q_unbuf <= my_rom(2414);
      when "100101101111" => q_unbuf <= my_rom(2415);
      when "100101110000" => q_unbuf <= my_rom(2416);
      when "100101110001" => q_unbuf <= my_rom(2417);
      when "100101110010" => q_unbuf <= my_rom(2418);
      when "100101110011" => q_unbuf <= my_rom(2419);
      when "100101110100" => q_unbuf <= my_rom(2420);
      when "100101110101" => q_unbuf <= my_rom(2421);
      when "100101110110" => q_unbuf <= my_rom(2422);
      when "100101110111" => q_unbuf <= my_rom(2423);
      when "100101111000" => q_unbuf <= my_rom(2424);
      when "100101111001" => q_unbuf <= my_rom(2425);
      when "100101111010" => q_unbuf <= my_rom(2426);
      when "100101111011" => q_unbuf <= my_rom(2427);
      when "100101111100" => q_unbuf <= my_rom(2428);
      when "100101111101" => q_unbuf <= my_rom(2429);
      when "100101111110" => q_unbuf <= my_rom(2430);
      when "100101111111" => q_unbuf <= my_rom(2431);
      when "100110000000" => q_unbuf <= my_rom(2432);
      when "100110000001" => q_unbuf <= my_rom(2433);
      when "100110000010" => q_unbuf <= my_rom(2434);
      when "100110000011" => q_unbuf <= my_rom(2435);
      when "100110000100" => q_unbuf <= my_rom(2436);
      when "100110000101" => q_unbuf <= my_rom(2437);
      when "100110000110" => q_unbuf <= my_rom(2438);
      when "100110000111" => q_unbuf <= my_rom(2439);
      when "100110001000" => q_unbuf <= my_rom(2440);
      when "100110001001" => q_unbuf <= my_rom(2441);
      when "100110001010" => q_unbuf <= my_rom(2442);
      when "100110001011" => q_unbuf <= my_rom(2443);
      when "100110001100" => q_unbuf <= my_rom(2444);
      when "100110001101" => q_unbuf <= my_rom(2445);
      when "100110001110" => q_unbuf <= my_rom(2446);
      when "100110001111" => q_unbuf <= my_rom(2447);
      when "100110010000" => q_unbuf <= my_rom(2448);
      when "100110010001" => q_unbuf <= my_rom(2449);
      when "100110010010" => q_unbuf <= my_rom(2450);
      when "100110010011" => q_unbuf <= my_rom(2451);
      when "100110010100" => q_unbuf <= my_rom(2452);
      when "100110010101" => q_unbuf <= my_rom(2453);
      when "100110010110" => q_unbuf <= my_rom(2454);
      when "100110010111" => q_unbuf <= my_rom(2455);
      when "100110011000" => q_unbuf <= my_rom(2456);
      when "100110011001" => q_unbuf <= my_rom(2457);
      when "100110011010" => q_unbuf <= my_rom(2458);
      when "100110011011" => q_unbuf <= my_rom(2459);
      when "100110011100" => q_unbuf <= my_rom(2460);
      when "100110011101" => q_unbuf <= my_rom(2461);
      when "100110011110" => q_unbuf <= my_rom(2462);
      when "100110011111" => q_unbuf <= my_rom(2463);
      when "100110100000" => q_unbuf <= my_rom(2464);
      when "100110100001" => q_unbuf <= my_rom(2465);
      when "100110100010" => q_unbuf <= my_rom(2466);
      when "100110100011" => q_unbuf <= my_rom(2467);
      when "100110100100" => q_unbuf <= my_rom(2468);
      when "100110100101" => q_unbuf <= my_rom(2469);
      when "100110100110" => q_unbuf <= my_rom(2470);
      when "100110100111" => q_unbuf <= my_rom(2471);
      when "100110101000" => q_unbuf <= my_rom(2472);
      when "100110101001" => q_unbuf <= my_rom(2473);
      when "100110101010" => q_unbuf <= my_rom(2474);
      when "100110101011" => q_unbuf <= my_rom(2475);
      when "100110101100" => q_unbuf <= my_rom(2476);
      when "100110101101" => q_unbuf <= my_rom(2477);
      when "100110101110" => q_unbuf <= my_rom(2478);
      when "100110101111" => q_unbuf <= my_rom(2479);
      when "100110110000" => q_unbuf <= my_rom(2480);
      when "100110110001" => q_unbuf <= my_rom(2481);
      when "100110110010" => q_unbuf <= my_rom(2482);
      when "100110110011" => q_unbuf <= my_rom(2483);
      when "100110110100" => q_unbuf <= my_rom(2484);
      when "100110110101" => q_unbuf <= my_rom(2485);
      when "100110110110" => q_unbuf <= my_rom(2486);
      when "100110110111" => q_unbuf <= my_rom(2487);
      when "100110111000" => q_unbuf <= my_rom(2488);
      when "100110111001" => q_unbuf <= my_rom(2489);
      when "100110111010" => q_unbuf <= my_rom(2490);
      when "100110111011" => q_unbuf <= my_rom(2491);
      when "100110111100" => q_unbuf <= my_rom(2492);
      when "100110111101" => q_unbuf <= my_rom(2493);
      when "100110111110" => q_unbuf <= my_rom(2494);
      when "100110111111" => q_unbuf <= my_rom(2495);
      when "100111000000" => q_unbuf <= my_rom(2496);
      when "100111000001" => q_unbuf <= my_rom(2497);
      when "100111000010" => q_unbuf <= my_rom(2498);
      when "100111000011" => q_unbuf <= my_rom(2499);
      when "100111000100" => q_unbuf <= my_rom(2500);
      when "100111000101" => q_unbuf <= my_rom(2501);
      when "100111000110" => q_unbuf <= my_rom(2502);
      when "100111000111" => q_unbuf <= my_rom(2503);
      when "100111001000" => q_unbuf <= my_rom(2504);
      when "100111001001" => q_unbuf <= my_rom(2505);
      when "100111001010" => q_unbuf <= my_rom(2506);
      when "100111001011" => q_unbuf <= my_rom(2507);
      when "100111001100" => q_unbuf <= my_rom(2508);
      when "100111001101" => q_unbuf <= my_rom(2509);
      when "100111001110" => q_unbuf <= my_rom(2510);
      when "100111001111" => q_unbuf <= my_rom(2511);
      when "100111010000" => q_unbuf <= my_rom(2512);
      when "100111010001" => q_unbuf <= my_rom(2513);
      when "100111010010" => q_unbuf <= my_rom(2514);
      when "100111010011" => q_unbuf <= my_rom(2515);
      when "100111010100" => q_unbuf <= my_rom(2516);
      when "100111010101" => q_unbuf <= my_rom(2517);
      when "100111010110" => q_unbuf <= my_rom(2518);
      when "100111010111" => q_unbuf <= my_rom(2519);
      when "100111011000" => q_unbuf <= my_rom(2520);
      when "100111011001" => q_unbuf <= my_rom(2521);
      when "100111011010" => q_unbuf <= my_rom(2522);
      when "100111011011" => q_unbuf <= my_rom(2523);
      when "100111011100" => q_unbuf <= my_rom(2524);
      when "100111011101" => q_unbuf <= my_rom(2525);
      when "100111011110" => q_unbuf <= my_rom(2526);
      when "100111011111" => q_unbuf <= my_rom(2527);
      when "100111100000" => q_unbuf <= my_rom(2528);
      when "100111100001" => q_unbuf <= my_rom(2529);
      when "100111100010" => q_unbuf <= my_rom(2530);
      when "100111100011" => q_unbuf <= my_rom(2531);
      when "100111100100" => q_unbuf <= my_rom(2532);
      when "100111100101" => q_unbuf <= my_rom(2533);
      when "100111100110" => q_unbuf <= my_rom(2534);
      when "100111100111" => q_unbuf <= my_rom(2535);
      when "100111101000" => q_unbuf <= my_rom(2536);
      when "100111101001" => q_unbuf <= my_rom(2537);
      when "100111101010" => q_unbuf <= my_rom(2538);
      when "100111101011" => q_unbuf <= my_rom(2539);
      when "100111101100" => q_unbuf <= my_rom(2540);
      when "100111101101" => q_unbuf <= my_rom(2541);
      when "100111101110" => q_unbuf <= my_rom(2542);
      when "100111101111" => q_unbuf <= my_rom(2543);
      when "100111110000" => q_unbuf <= my_rom(2544);
      when "100111110001" => q_unbuf <= my_rom(2545);
      when "100111110010" => q_unbuf <= my_rom(2546);
      when "100111110011" => q_unbuf <= my_rom(2547);
      when "100111110100" => q_unbuf <= my_rom(2548);
      when "100111110101" => q_unbuf <= my_rom(2549);
      when "100111110110" => q_unbuf <= my_rom(2550);
      when "100111110111" => q_unbuf <= my_rom(2551);
      when "100111111000" => q_unbuf <= my_rom(2552);
      when "100111111001" => q_unbuf <= my_rom(2553);
      when "100111111010" => q_unbuf <= my_rom(2554);
      when "100111111011" => q_unbuf <= my_rom(2555);
      when "100111111100" => q_unbuf <= my_rom(2556);
      when "100111111101" => q_unbuf <= my_rom(2557);
      when "100111111110" => q_unbuf <= my_rom(2558);
      when "100111111111" => q_unbuf <= my_rom(2559);
      when "101000000000" => q_unbuf <= my_rom(2560);
      when "101000000001" => q_unbuf <= my_rom(2561);
      when "101000000010" => q_unbuf <= my_rom(2562);
      when "101000000011" => q_unbuf <= my_rom(2563);
      when "101000000100" => q_unbuf <= my_rom(2564);
      when "101000000101" => q_unbuf <= my_rom(2565);
      when "101000000110" => q_unbuf <= my_rom(2566);
      when "101000000111" => q_unbuf <= my_rom(2567);
      when "101000001000" => q_unbuf <= my_rom(2568);
      when "101000001001" => q_unbuf <= my_rom(2569);
      when "101000001010" => q_unbuf <= my_rom(2570);
      when "101000001011" => q_unbuf <= my_rom(2571);
      when "101000001100" => q_unbuf <= my_rom(2572);
      when "101000001101" => q_unbuf <= my_rom(2573);
      when "101000001110" => q_unbuf <= my_rom(2574);
      when "101000001111" => q_unbuf <= my_rom(2575);
      when "101000010000" => q_unbuf <= my_rom(2576);
      when "101000010001" => q_unbuf <= my_rom(2577);
      when "101000010010" => q_unbuf <= my_rom(2578);
      when "101000010011" => q_unbuf <= my_rom(2579);
      when "101000010100" => q_unbuf <= my_rom(2580);
      when "101000010101" => q_unbuf <= my_rom(2581);
      when "101000010110" => q_unbuf <= my_rom(2582);
      when "101000010111" => q_unbuf <= my_rom(2583);
      when "101000011000" => q_unbuf <= my_rom(2584);
      when "101000011001" => q_unbuf <= my_rom(2585);
      when "101000011010" => q_unbuf <= my_rom(2586);
      when "101000011011" => q_unbuf <= my_rom(2587);
      when "101000011100" => q_unbuf <= my_rom(2588);
      when "101000011101" => q_unbuf <= my_rom(2589);
      when "101000011110" => q_unbuf <= my_rom(2590);
      when "101000011111" => q_unbuf <= my_rom(2591);
      when "101000100000" => q_unbuf <= my_rom(2592);
      when "101000100001" => q_unbuf <= my_rom(2593);
      when "101000100010" => q_unbuf <= my_rom(2594);
      when "101000100011" => q_unbuf <= my_rom(2595);
      when "101000100100" => q_unbuf <= my_rom(2596);
      when "101000100101" => q_unbuf <= my_rom(2597);
      when "101000100110" => q_unbuf <= my_rom(2598);
      when "101000100111" => q_unbuf <= my_rom(2599);
      when "101000101000" => q_unbuf <= my_rom(2600);
      when "101000101001" => q_unbuf <= my_rom(2601);
      when "101000101010" => q_unbuf <= my_rom(2602);
      when "101000101011" => q_unbuf <= my_rom(2603);
      when "101000101100" => q_unbuf <= my_rom(2604);
      when "101000101101" => q_unbuf <= my_rom(2605);
      when "101000101110" => q_unbuf <= my_rom(2606);
      when "101000101111" => q_unbuf <= my_rom(2607);
      when "101000110000" => q_unbuf <= my_rom(2608);
      when "101000110001" => q_unbuf <= my_rom(2609);
      when "101000110010" => q_unbuf <= my_rom(2610);
      when "101000110011" => q_unbuf <= my_rom(2611);
      when "101000110100" => q_unbuf <= my_rom(2612);
      when "101000110101" => q_unbuf <= my_rom(2613);
      when "101000110110" => q_unbuf <= my_rom(2614);
      when "101000110111" => q_unbuf <= my_rom(2615);
      when "101000111000" => q_unbuf <= my_rom(2616);
      when "101000111001" => q_unbuf <= my_rom(2617);
      when "101000111010" => q_unbuf <= my_rom(2618);
      when "101000111011" => q_unbuf <= my_rom(2619);
      when "101000111100" => q_unbuf <= my_rom(2620);
      when "101000111101" => q_unbuf <= my_rom(2621);
      when "101000111110" => q_unbuf <= my_rom(2622);
      when "101000111111" => q_unbuf <= my_rom(2623);
      when "101001000000" => q_unbuf <= my_rom(2624);
      when "101001000001" => q_unbuf <= my_rom(2625);
      when "101001000010" => q_unbuf <= my_rom(2626);
      when "101001000011" => q_unbuf <= my_rom(2627);
      when "101001000100" => q_unbuf <= my_rom(2628);
      when "101001000101" => q_unbuf <= my_rom(2629);
      when "101001000110" => q_unbuf <= my_rom(2630);
      when "101001000111" => q_unbuf <= my_rom(2631);
      when "101001001000" => q_unbuf <= my_rom(2632);
      when "101001001001" => q_unbuf <= my_rom(2633);
      when "101001001010" => q_unbuf <= my_rom(2634);
      when "101001001011" => q_unbuf <= my_rom(2635);
      when "101001001100" => q_unbuf <= my_rom(2636);
      when "101001001101" => q_unbuf <= my_rom(2637);
      when "101001001110" => q_unbuf <= my_rom(2638);
      when "101001001111" => q_unbuf <= my_rom(2639);
      when "101001010000" => q_unbuf <= my_rom(2640);
      when "101001010001" => q_unbuf <= my_rom(2641);
      when "101001010010" => q_unbuf <= my_rom(2642);
      when "101001010011" => q_unbuf <= my_rom(2643);
      when "101001010100" => q_unbuf <= my_rom(2644);
      when "101001010101" => q_unbuf <= my_rom(2645);
      when "101001010110" => q_unbuf <= my_rom(2646);
      when "101001010111" => q_unbuf <= my_rom(2647);
      when "101001011000" => q_unbuf <= my_rom(2648);
      when "101001011001" => q_unbuf <= my_rom(2649);
      when "101001011010" => q_unbuf <= my_rom(2650);
      when "101001011011" => q_unbuf <= my_rom(2651);
      when "101001011100" => q_unbuf <= my_rom(2652);
      when "101001011101" => q_unbuf <= my_rom(2653);
      when "101001011110" => q_unbuf <= my_rom(2654);
      when "101001011111" => q_unbuf <= my_rom(2655);
      when "101001100000" => q_unbuf <= my_rom(2656);
      when "101001100001" => q_unbuf <= my_rom(2657);
      when "101001100010" => q_unbuf <= my_rom(2658);
      when "101001100011" => q_unbuf <= my_rom(2659);
      when "101001100100" => q_unbuf <= my_rom(2660);
      when "101001100101" => q_unbuf <= my_rom(2661);
      when "101001100110" => q_unbuf <= my_rom(2662);
      when "101001100111" => q_unbuf <= my_rom(2663);
      when "101001101000" => q_unbuf <= my_rom(2664);
      when "101001101001" => q_unbuf <= my_rom(2665);
      when "101001101010" => q_unbuf <= my_rom(2666);
      when "101001101011" => q_unbuf <= my_rom(2667);
      when "101001101100" => q_unbuf <= my_rom(2668);
      when "101001101101" => q_unbuf <= my_rom(2669);
      when "101001101110" => q_unbuf <= my_rom(2670);
      when "101001101111" => q_unbuf <= my_rom(2671);
      when "101001110000" => q_unbuf <= my_rom(2672);
      when "101001110001" => q_unbuf <= my_rom(2673);
      when "101001110010" => q_unbuf <= my_rom(2674);
      when "101001110011" => q_unbuf <= my_rom(2675);
      when "101001110100" => q_unbuf <= my_rom(2676);
      when "101001110101" => q_unbuf <= my_rom(2677);
      when "101001110110" => q_unbuf <= my_rom(2678);
      when "101001110111" => q_unbuf <= my_rom(2679);
      when "101001111000" => q_unbuf <= my_rom(2680);
      when "101001111001" => q_unbuf <= my_rom(2681);
      when "101001111010" => q_unbuf <= my_rom(2682);
      when "101001111011" => q_unbuf <= my_rom(2683);
      when "101001111100" => q_unbuf <= my_rom(2684);
      when "101001111101" => q_unbuf <= my_rom(2685);
      when "101001111110" => q_unbuf <= my_rom(2686);
      when "101001111111" => q_unbuf <= my_rom(2687);
      when "101010000000" => q_unbuf <= my_rom(2688);
      when "101010000001" => q_unbuf <= my_rom(2689);
      when "101010000010" => q_unbuf <= my_rom(2690);
      when "101010000011" => q_unbuf <= my_rom(2691);
      when "101010000100" => q_unbuf <= my_rom(2692);
      when "101010000101" => q_unbuf <= my_rom(2693);
      when "101010000110" => q_unbuf <= my_rom(2694);
      when "101010000111" => q_unbuf <= my_rom(2695);
      when "101010001000" => q_unbuf <= my_rom(2696);
      when "101010001001" => q_unbuf <= my_rom(2697);
      when "101010001010" => q_unbuf <= my_rom(2698);
      when "101010001011" => q_unbuf <= my_rom(2699);
      when "101010001100" => q_unbuf <= my_rom(2700);
      when "101010001101" => q_unbuf <= my_rom(2701);
      when "101010001110" => q_unbuf <= my_rom(2702);
      when "101010001111" => q_unbuf <= my_rom(2703);
      when "101010010000" => q_unbuf <= my_rom(2704);
      when "101010010001" => q_unbuf <= my_rom(2705);
      when "101010010010" => q_unbuf <= my_rom(2706);
      when "101010010011" => q_unbuf <= my_rom(2707);
      when "101010010100" => q_unbuf <= my_rom(2708);
      when "101010010101" => q_unbuf <= my_rom(2709);
      when "101010010110" => q_unbuf <= my_rom(2710);
      when "101010010111" => q_unbuf <= my_rom(2711);
      when "101010011000" => q_unbuf <= my_rom(2712);
      when "101010011001" => q_unbuf <= my_rom(2713);
      when "101010011010" => q_unbuf <= my_rom(2714);
      when "101010011011" => q_unbuf <= my_rom(2715);
      when "101010011100" => q_unbuf <= my_rom(2716);
      when "101010011101" => q_unbuf <= my_rom(2717);
      when "101010011110" => q_unbuf <= my_rom(2718);
      when "101010011111" => q_unbuf <= my_rom(2719);
      when "101010100000" => q_unbuf <= my_rom(2720);
      when "101010100001" => q_unbuf <= my_rom(2721);
      when "101010100010" => q_unbuf <= my_rom(2722);
      when "101010100011" => q_unbuf <= my_rom(2723);
      when "101010100100" => q_unbuf <= my_rom(2724);
      when "101010100101" => q_unbuf <= my_rom(2725);
      when "101010100110" => q_unbuf <= my_rom(2726);
      when "101010100111" => q_unbuf <= my_rom(2727);
      when "101010101000" => q_unbuf <= my_rom(2728);
      when "101010101001" => q_unbuf <= my_rom(2729);
      when "101010101010" => q_unbuf <= my_rom(2730);
      when "101010101011" => q_unbuf <= my_rom(2731);
      when "101010101100" => q_unbuf <= my_rom(2732);
      when "101010101101" => q_unbuf <= my_rom(2733);
      when "101010101110" => q_unbuf <= my_rom(2734);
      when "101010101111" => q_unbuf <= my_rom(2735);
      when "101010110000" => q_unbuf <= my_rom(2736);
      when "101010110001" => q_unbuf <= my_rom(2737);
      when "101010110010" => q_unbuf <= my_rom(2738);
      when "101010110011" => q_unbuf <= my_rom(2739);
      when "101010110100" => q_unbuf <= my_rom(2740);
      when "101010110101" => q_unbuf <= my_rom(2741);
      when "101010110110" => q_unbuf <= my_rom(2742);
      when "101010110111" => q_unbuf <= my_rom(2743);
      when "101010111000" => q_unbuf <= my_rom(2744);
      when "101010111001" => q_unbuf <= my_rom(2745);
      when "101010111010" => q_unbuf <= my_rom(2746);
      when "101010111011" => q_unbuf <= my_rom(2747);
      when "101010111100" => q_unbuf <= my_rom(2748);
      when "101010111101" => q_unbuf <= my_rom(2749);
      when "101010111110" => q_unbuf <= my_rom(2750);
      when "101010111111" => q_unbuf <= my_rom(2751);
      when "101011000000" => q_unbuf <= my_rom(2752);
      when "101011000001" => q_unbuf <= my_rom(2753);
      when "101011000010" => q_unbuf <= my_rom(2754);
      when "101011000011" => q_unbuf <= my_rom(2755);
      when "101011000100" => q_unbuf <= my_rom(2756);
      when "101011000101" => q_unbuf <= my_rom(2757);
      when "101011000110" => q_unbuf <= my_rom(2758);
      when "101011000111" => q_unbuf <= my_rom(2759);
      when "101011001000" => q_unbuf <= my_rom(2760);
      when "101011001001" => q_unbuf <= my_rom(2761);
      when "101011001010" => q_unbuf <= my_rom(2762);
      when "101011001011" => q_unbuf <= my_rom(2763);
      when "101011001100" => q_unbuf <= my_rom(2764);
      when "101011001101" => q_unbuf <= my_rom(2765);
      when "101011001110" => q_unbuf <= my_rom(2766);
      when "101011001111" => q_unbuf <= my_rom(2767);
      when "101011010000" => q_unbuf <= my_rom(2768);
      when "101011010001" => q_unbuf <= my_rom(2769);
      when "101011010010" => q_unbuf <= my_rom(2770);
      when "101011010011" => q_unbuf <= my_rom(2771);
      when "101011010100" => q_unbuf <= my_rom(2772);
      when "101011010101" => q_unbuf <= my_rom(2773);
      when "101011010110" => q_unbuf <= my_rom(2774);
      when "101011010111" => q_unbuf <= my_rom(2775);
      when "101011011000" => q_unbuf <= my_rom(2776);
      when "101011011001" => q_unbuf <= my_rom(2777);
      when "101011011010" => q_unbuf <= my_rom(2778);
      when "101011011011" => q_unbuf <= my_rom(2779);
      when "101011011100" => q_unbuf <= my_rom(2780);
      when "101011011101" => q_unbuf <= my_rom(2781);
      when "101011011110" => q_unbuf <= my_rom(2782);
      when "101011011111" => q_unbuf <= my_rom(2783);
      when "101011100000" => q_unbuf <= my_rom(2784);
      when "101011100001" => q_unbuf <= my_rom(2785);
      when "101011100010" => q_unbuf <= my_rom(2786);
      when "101011100011" => q_unbuf <= my_rom(2787);
      when "101011100100" => q_unbuf <= my_rom(2788);
      when "101011100101" => q_unbuf <= my_rom(2789);
      when "101011100110" => q_unbuf <= my_rom(2790);
      when "101011100111" => q_unbuf <= my_rom(2791);
      when "101011101000" => q_unbuf <= my_rom(2792);
      when "101011101001" => q_unbuf <= my_rom(2793);
      when "101011101010" => q_unbuf <= my_rom(2794);
      when "101011101011" => q_unbuf <= my_rom(2795);
      when "101011101100" => q_unbuf <= my_rom(2796);
      when "101011101101" => q_unbuf <= my_rom(2797);
      when "101011101110" => q_unbuf <= my_rom(2798);
      when "101011101111" => q_unbuf <= my_rom(2799);
      when "101011110000" => q_unbuf <= my_rom(2800);
      when "101011110001" => q_unbuf <= my_rom(2801);
      when "101011110010" => q_unbuf <= my_rom(2802);
      when "101011110011" => q_unbuf <= my_rom(2803);
      when "101011110100" => q_unbuf <= my_rom(2804);
      when "101011110101" => q_unbuf <= my_rom(2805);
      when "101011110110" => q_unbuf <= my_rom(2806);
      when "101011110111" => q_unbuf <= my_rom(2807);
      when "101011111000" => q_unbuf <= my_rom(2808);
      when "101011111001" => q_unbuf <= my_rom(2809);
      when "101011111010" => q_unbuf <= my_rom(2810);
      when "101011111011" => q_unbuf <= my_rom(2811);
      when "101011111100" => q_unbuf <= my_rom(2812);
      when "101011111101" => q_unbuf <= my_rom(2813);
      when "101011111110" => q_unbuf <= my_rom(2814);
      when "101011111111" => q_unbuf <= my_rom(2815);
      when "101100000000" => q_unbuf <= my_rom(2816);
      when "101100000001" => q_unbuf <= my_rom(2817);
      when "101100000010" => q_unbuf <= my_rom(2818);
      when "101100000011" => q_unbuf <= my_rom(2819);
      when "101100000100" => q_unbuf <= my_rom(2820);
      when "101100000101" => q_unbuf <= my_rom(2821);
      when "101100000110" => q_unbuf <= my_rom(2822);
      when "101100000111" => q_unbuf <= my_rom(2823);
      when "101100001000" => q_unbuf <= my_rom(2824);
      when "101100001001" => q_unbuf <= my_rom(2825);
      when "101100001010" => q_unbuf <= my_rom(2826);
      when "101100001011" => q_unbuf <= my_rom(2827);
      when "101100001100" => q_unbuf <= my_rom(2828);
      when "101100001101" => q_unbuf <= my_rom(2829);
      when "101100001110" => q_unbuf <= my_rom(2830);
      when "101100001111" => q_unbuf <= my_rom(2831);
      when "101100010000" => q_unbuf <= my_rom(2832);
      when "101100010001" => q_unbuf <= my_rom(2833);
      when "101100010010" => q_unbuf <= my_rom(2834);
      when "101100010011" => q_unbuf <= my_rom(2835);
      when "101100010100" => q_unbuf <= my_rom(2836);
      when "101100010101" => q_unbuf <= my_rom(2837);
      when "101100010110" => q_unbuf <= my_rom(2838);
      when "101100010111" => q_unbuf <= my_rom(2839);
      when "101100011000" => q_unbuf <= my_rom(2840);
      when "101100011001" => q_unbuf <= my_rom(2841);
      when "101100011010" => q_unbuf <= my_rom(2842);
      when "101100011011" => q_unbuf <= my_rom(2843);
      when "101100011100" => q_unbuf <= my_rom(2844);
      when "101100011101" => q_unbuf <= my_rom(2845);
      when "101100011110" => q_unbuf <= my_rom(2846);
      when "101100011111" => q_unbuf <= my_rom(2847);
      when "101100100000" => q_unbuf <= my_rom(2848);
      when "101100100001" => q_unbuf <= my_rom(2849);
      when "101100100010" => q_unbuf <= my_rom(2850);
      when "101100100011" => q_unbuf <= my_rom(2851);
      when "101100100100" => q_unbuf <= my_rom(2852);
      when "101100100101" => q_unbuf <= my_rom(2853);
      when "101100100110" => q_unbuf <= my_rom(2854);
      when "101100100111" => q_unbuf <= my_rom(2855);
      when "101100101000" => q_unbuf <= my_rom(2856);
      when "101100101001" => q_unbuf <= my_rom(2857);
      when "101100101010" => q_unbuf <= my_rom(2858);
      when "101100101011" => q_unbuf <= my_rom(2859);
      when "101100101100" => q_unbuf <= my_rom(2860);
      when "101100101101" => q_unbuf <= my_rom(2861);
      when "101100101110" => q_unbuf <= my_rom(2862);
      when "101100101111" => q_unbuf <= my_rom(2863);
      when "101100110000" => q_unbuf <= my_rom(2864);
      when "101100110001" => q_unbuf <= my_rom(2865);
      when "101100110010" => q_unbuf <= my_rom(2866);
      when "101100110011" => q_unbuf <= my_rom(2867);
      when "101100110100" => q_unbuf <= my_rom(2868);
      when "101100110101" => q_unbuf <= my_rom(2869);
      when "101100110110" => q_unbuf <= my_rom(2870);
      when "101100110111" => q_unbuf <= my_rom(2871);
      when "101100111000" => q_unbuf <= my_rom(2872);
      when "101100111001" => q_unbuf <= my_rom(2873);
      when "101100111010" => q_unbuf <= my_rom(2874);
      when "101100111011" => q_unbuf <= my_rom(2875);
      when "101100111100" => q_unbuf <= my_rom(2876);
      when "101100111101" => q_unbuf <= my_rom(2877);
      when "101100111110" => q_unbuf <= my_rom(2878);
      when "101100111111" => q_unbuf <= my_rom(2879);
      when "101101000000" => q_unbuf <= my_rom(2880);
      when "101101000001" => q_unbuf <= my_rom(2881);
      when "101101000010" => q_unbuf <= my_rom(2882);
      when "101101000011" => q_unbuf <= my_rom(2883);
      when "101101000100" => q_unbuf <= my_rom(2884);
      when "101101000101" => q_unbuf <= my_rom(2885);
      when "101101000110" => q_unbuf <= my_rom(2886);
      when "101101000111" => q_unbuf <= my_rom(2887);
      when "101101001000" => q_unbuf <= my_rom(2888);
      when "101101001001" => q_unbuf <= my_rom(2889);
      when "101101001010" => q_unbuf <= my_rom(2890);
      when "101101001011" => q_unbuf <= my_rom(2891);
      when "101101001100" => q_unbuf <= my_rom(2892);
      when "101101001101" => q_unbuf <= my_rom(2893);
      when "101101001110" => q_unbuf <= my_rom(2894);
      when "101101001111" => q_unbuf <= my_rom(2895);
      when "101101010000" => q_unbuf <= my_rom(2896);
      when "101101010001" => q_unbuf <= my_rom(2897);
      when "101101010010" => q_unbuf <= my_rom(2898);
      when "101101010011" => q_unbuf <= my_rom(2899);
      when "101101010100" => q_unbuf <= my_rom(2900);
      when "101101010101" => q_unbuf <= my_rom(2901);
      when "101101010110" => q_unbuf <= my_rom(2902);
      when "101101010111" => q_unbuf <= my_rom(2903);
      when "101101011000" => q_unbuf <= my_rom(2904);
      when "101101011001" => q_unbuf <= my_rom(2905);
      when "101101011010" => q_unbuf <= my_rom(2906);
      when "101101011011" => q_unbuf <= my_rom(2907);
      when "101101011100" => q_unbuf <= my_rom(2908);
      when "101101011101" => q_unbuf <= my_rom(2909);
      when "101101011110" => q_unbuf <= my_rom(2910);
      when "101101011111" => q_unbuf <= my_rom(2911);
      when "101101100000" => q_unbuf <= my_rom(2912);
      when "101101100001" => q_unbuf <= my_rom(2913);
      when "101101100010" => q_unbuf <= my_rom(2914);
      when "101101100011" => q_unbuf <= my_rom(2915);
      when "101101100100" => q_unbuf <= my_rom(2916);
      when "101101100101" => q_unbuf <= my_rom(2917);
      when "101101100110" => q_unbuf <= my_rom(2918);
      when "101101100111" => q_unbuf <= my_rom(2919);
      when "101101101000" => q_unbuf <= my_rom(2920);
      when "101101101001" => q_unbuf <= my_rom(2921);
      when "101101101010" => q_unbuf <= my_rom(2922);
      when "101101101011" => q_unbuf <= my_rom(2923);
      when "101101101100" => q_unbuf <= my_rom(2924);
      when "101101101101" => q_unbuf <= my_rom(2925);
      when "101101101110" => q_unbuf <= my_rom(2926);
      when "101101101111" => q_unbuf <= my_rom(2927);
      when "101101110000" => q_unbuf <= my_rom(2928);
      when "101101110001" => q_unbuf <= my_rom(2929);
      when "101101110010" => q_unbuf <= my_rom(2930);
      when "101101110011" => q_unbuf <= my_rom(2931);
      when "101101110100" => q_unbuf <= my_rom(2932);
      when "101101110101" => q_unbuf <= my_rom(2933);
      when "101101110110" => q_unbuf <= my_rom(2934);
      when "101101110111" => q_unbuf <= my_rom(2935);
      when "101101111000" => q_unbuf <= my_rom(2936);
      when "101101111001" => q_unbuf <= my_rom(2937);
      when "101101111010" => q_unbuf <= my_rom(2938);
      when "101101111011" => q_unbuf <= my_rom(2939);
      when "101101111100" => q_unbuf <= my_rom(2940);
      when "101101111101" => q_unbuf <= my_rom(2941);
      when "101101111110" => q_unbuf <= my_rom(2942);
      when "101101111111" => q_unbuf <= my_rom(2943);
      when "101110000000" => q_unbuf <= my_rom(2944);
      when "101110000001" => q_unbuf <= my_rom(2945);
      when "101110000010" => q_unbuf <= my_rom(2946);
      when "101110000011" => q_unbuf <= my_rom(2947);
      when "101110000100" => q_unbuf <= my_rom(2948);
      when "101110000101" => q_unbuf <= my_rom(2949);
      when "101110000110" => q_unbuf <= my_rom(2950);
      when "101110000111" => q_unbuf <= my_rom(2951);
      when "101110001000" => q_unbuf <= my_rom(2952);
      when "101110001001" => q_unbuf <= my_rom(2953);
      when "101110001010" => q_unbuf <= my_rom(2954);
      when "101110001011" => q_unbuf <= my_rom(2955);
      when "101110001100" => q_unbuf <= my_rom(2956);
      when "101110001101" => q_unbuf <= my_rom(2957);
      when "101110001110" => q_unbuf <= my_rom(2958);
      when "101110001111" => q_unbuf <= my_rom(2959);
      when "101110010000" => q_unbuf <= my_rom(2960);
      when "101110010001" => q_unbuf <= my_rom(2961);
      when "101110010010" => q_unbuf <= my_rom(2962);
      when "101110010011" => q_unbuf <= my_rom(2963);
      when "101110010100" => q_unbuf <= my_rom(2964);
      when "101110010101" => q_unbuf <= my_rom(2965);
      when "101110010110" => q_unbuf <= my_rom(2966);
      when "101110010111" => q_unbuf <= my_rom(2967);
      when "101110011000" => q_unbuf <= my_rom(2968);
      when "101110011001" => q_unbuf <= my_rom(2969);
      when "101110011010" => q_unbuf <= my_rom(2970);
      when "101110011011" => q_unbuf <= my_rom(2971);
      when "101110011100" => q_unbuf <= my_rom(2972);
      when "101110011101" => q_unbuf <= my_rom(2973);
      when "101110011110" => q_unbuf <= my_rom(2974);
      when "101110011111" => q_unbuf <= my_rom(2975);
      when "101110100000" => q_unbuf <= my_rom(2976);
      when "101110100001" => q_unbuf <= my_rom(2977);
      when "101110100010" => q_unbuf <= my_rom(2978);
      when "101110100011" => q_unbuf <= my_rom(2979);
      when "101110100100" => q_unbuf <= my_rom(2980);
      when "101110100101" => q_unbuf <= my_rom(2981);
      when "101110100110" => q_unbuf <= my_rom(2982);
      when "101110100111" => q_unbuf <= my_rom(2983);
      when "101110101000" => q_unbuf <= my_rom(2984);
      when "101110101001" => q_unbuf <= my_rom(2985);
      when "101110101010" => q_unbuf <= my_rom(2986);
      when "101110101011" => q_unbuf <= my_rom(2987);
      when "101110101100" => q_unbuf <= my_rom(2988);
      when "101110101101" => q_unbuf <= my_rom(2989);
      when "101110101110" => q_unbuf <= my_rom(2990);
      when "101110101111" => q_unbuf <= my_rom(2991);
      when "101110110000" => q_unbuf <= my_rom(2992);
      when "101110110001" => q_unbuf <= my_rom(2993);
      when "101110110010" => q_unbuf <= my_rom(2994);
      when "101110110011" => q_unbuf <= my_rom(2995);
      when "101110110100" => q_unbuf <= my_rom(2996);
      when "101110110101" => q_unbuf <= my_rom(2997);
      when "101110110110" => q_unbuf <= my_rom(2998);
      when "101110110111" => q_unbuf <= my_rom(2999);
      when "101110111000" => q_unbuf <= my_rom(3000);
      when "101110111001" => q_unbuf <= my_rom(3001);
      when "101110111010" => q_unbuf <= my_rom(3002);
      when "101110111011" => q_unbuf <= my_rom(3003);
      when "101110111100" => q_unbuf <= my_rom(3004);
      when "101110111101" => q_unbuf <= my_rom(3005);
      when "101110111110" => q_unbuf <= my_rom(3006);
      when "101110111111" => q_unbuf <= my_rom(3007);
      when "101111000000" => q_unbuf <= my_rom(3008);
      when "101111000001" => q_unbuf <= my_rom(3009);
      when "101111000010" => q_unbuf <= my_rom(3010);
      when "101111000011" => q_unbuf <= my_rom(3011);
      when "101111000100" => q_unbuf <= my_rom(3012);
      when "101111000101" => q_unbuf <= my_rom(3013);
      when "101111000110" => q_unbuf <= my_rom(3014);
      when "101111000111" => q_unbuf <= my_rom(3015);
      when "101111001000" => q_unbuf <= my_rom(3016);
      when "101111001001" => q_unbuf <= my_rom(3017);
      when "101111001010" => q_unbuf <= my_rom(3018);
      when "101111001011" => q_unbuf <= my_rom(3019);
      when "101111001100" => q_unbuf <= my_rom(3020);
      when "101111001101" => q_unbuf <= my_rom(3021);
      when "101111001110" => q_unbuf <= my_rom(3022);
      when "101111001111" => q_unbuf <= my_rom(3023);
      when "101111010000" => q_unbuf <= my_rom(3024);
      when "101111010001" => q_unbuf <= my_rom(3025);
      when "101111010010" => q_unbuf <= my_rom(3026);
      when "101111010011" => q_unbuf <= my_rom(3027);
      when "101111010100" => q_unbuf <= my_rom(3028);
      when "101111010101" => q_unbuf <= my_rom(3029);
      when "101111010110" => q_unbuf <= my_rom(3030);
      when "101111010111" => q_unbuf <= my_rom(3031);
      when "101111011000" => q_unbuf <= my_rom(3032);
      when "101111011001" => q_unbuf <= my_rom(3033);
      when "101111011010" => q_unbuf <= my_rom(3034);
      when "101111011011" => q_unbuf <= my_rom(3035);
      when "101111011100" => q_unbuf <= my_rom(3036);
      when "101111011101" => q_unbuf <= my_rom(3037);
      when "101111011110" => q_unbuf <= my_rom(3038);
      when "101111011111" => q_unbuf <= my_rom(3039);
      when "101111100000" => q_unbuf <= my_rom(3040);
      when "101111100001" => q_unbuf <= my_rom(3041);
      when "101111100010" => q_unbuf <= my_rom(3042);
      when "101111100011" => q_unbuf <= my_rom(3043);
      when "101111100100" => q_unbuf <= my_rom(3044);
      when "101111100101" => q_unbuf <= my_rom(3045);
      when "101111100110" => q_unbuf <= my_rom(3046);
      when "101111100111" => q_unbuf <= my_rom(3047);
      when "101111101000" => q_unbuf <= my_rom(3048);
      when "101111101001" => q_unbuf <= my_rom(3049);
      when "101111101010" => q_unbuf <= my_rom(3050);
      when "101111101011" => q_unbuf <= my_rom(3051);
      when "101111101100" => q_unbuf <= my_rom(3052);
      when "101111101101" => q_unbuf <= my_rom(3053);
      when "101111101110" => q_unbuf <= my_rom(3054);
      when "101111101111" => q_unbuf <= my_rom(3055);
      when "101111110000" => q_unbuf <= my_rom(3056);
      when "101111110001" => q_unbuf <= my_rom(3057);
      when "101111110010" => q_unbuf <= my_rom(3058);
      when "101111110011" => q_unbuf <= my_rom(3059);
      when "101111110100" => q_unbuf <= my_rom(3060);
      when "101111110101" => q_unbuf <= my_rom(3061);
      when "101111110110" => q_unbuf <= my_rom(3062);
      when "101111110111" => q_unbuf <= my_rom(3063);
      when "101111111000" => q_unbuf <= my_rom(3064);
      when "101111111001" => q_unbuf <= my_rom(3065);
      when "101111111010" => q_unbuf <= my_rom(3066);
      when "101111111011" => q_unbuf <= my_rom(3067);
      when "101111111100" => q_unbuf <= my_rom(3068);
      when "101111111101" => q_unbuf <= my_rom(3069);
      when "101111111110" => q_unbuf <= my_rom(3070);
      when "101111111111" => q_unbuf <= my_rom(3071);
      when "110000000000" => q_unbuf <= my_rom(3072);
      when "110000000001" => q_unbuf <= my_rom(3073);
      when "110000000010" => q_unbuf <= my_rom(3074);
      when "110000000011" => q_unbuf <= my_rom(3075);
      when "110000000100" => q_unbuf <= my_rom(3076);
      when "110000000101" => q_unbuf <= my_rom(3077);
      when "110000000110" => q_unbuf <= my_rom(3078);
      when "110000000111" => q_unbuf <= my_rom(3079);
      when "110000001000" => q_unbuf <= my_rom(3080);
      when "110000001001" => q_unbuf <= my_rom(3081);
      when "110000001010" => q_unbuf <= my_rom(3082);
      when "110000001011" => q_unbuf <= my_rom(3083);
      when "110000001100" => q_unbuf <= my_rom(3084);
      when "110000001101" => q_unbuf <= my_rom(3085);
      when "110000001110" => q_unbuf <= my_rom(3086);
      when "110000001111" => q_unbuf <= my_rom(3087);
      when "110000010000" => q_unbuf <= my_rom(3088);
      when "110000010001" => q_unbuf <= my_rom(3089);
      when "110000010010" => q_unbuf <= my_rom(3090);
      when "110000010011" => q_unbuf <= my_rom(3091);
      when "110000010100" => q_unbuf <= my_rom(3092);
      when "110000010101" => q_unbuf <= my_rom(3093);
      when "110000010110" => q_unbuf <= my_rom(3094);
      when "110000010111" => q_unbuf <= my_rom(3095);
      when "110000011000" => q_unbuf <= my_rom(3096);
      when "110000011001" => q_unbuf <= my_rom(3097);
      when "110000011010" => q_unbuf <= my_rom(3098);
      when "110000011011" => q_unbuf <= my_rom(3099);
      when "110000011100" => q_unbuf <= my_rom(3100);
      when "110000011101" => q_unbuf <= my_rom(3101);
      when "110000011110" => q_unbuf <= my_rom(3102);
      when "110000011111" => q_unbuf <= my_rom(3103);
      when "110000100000" => q_unbuf <= my_rom(3104);
      when "110000100001" => q_unbuf <= my_rom(3105);
      when "110000100010" => q_unbuf <= my_rom(3106);
      when "110000100011" => q_unbuf <= my_rom(3107);
      when "110000100100" => q_unbuf <= my_rom(3108);
      when "110000100101" => q_unbuf <= my_rom(3109);
      when "110000100110" => q_unbuf <= my_rom(3110);
      when "110000100111" => q_unbuf <= my_rom(3111);
      when "110000101000" => q_unbuf <= my_rom(3112);
      when "110000101001" => q_unbuf <= my_rom(3113);
      when "110000101010" => q_unbuf <= my_rom(3114);
      when "110000101011" => q_unbuf <= my_rom(3115);
      when "110000101100" => q_unbuf <= my_rom(3116);
      when "110000101101" => q_unbuf <= my_rom(3117);
      when "110000101110" => q_unbuf <= my_rom(3118);
      when "110000101111" => q_unbuf <= my_rom(3119);
      when "110000110000" => q_unbuf <= my_rom(3120);
      when "110000110001" => q_unbuf <= my_rom(3121);
      when "110000110010" => q_unbuf <= my_rom(3122);
      when "110000110011" => q_unbuf <= my_rom(3123);
      when "110000110100" => q_unbuf <= my_rom(3124);
      when "110000110101" => q_unbuf <= my_rom(3125);
      when "110000110110" => q_unbuf <= my_rom(3126);
      when "110000110111" => q_unbuf <= my_rom(3127);
      when "110000111000" => q_unbuf <= my_rom(3128);
      when "110000111001" => q_unbuf <= my_rom(3129);
      when "110000111010" => q_unbuf <= my_rom(3130);
      when "110000111011" => q_unbuf <= my_rom(3131);
      when "110000111100" => q_unbuf <= my_rom(3132);
      when "110000111101" => q_unbuf <= my_rom(3133);
      when "110000111110" => q_unbuf <= my_rom(3134);
      when "110000111111" => q_unbuf <= my_rom(3135);
      when "110001000000" => q_unbuf <= my_rom(3136);
      when "110001000001" => q_unbuf <= my_rom(3137);
      when "110001000010" => q_unbuf <= my_rom(3138);
      when "110001000011" => q_unbuf <= my_rom(3139);
      when "110001000100" => q_unbuf <= my_rom(3140);
      when "110001000101" => q_unbuf <= my_rom(3141);
      when "110001000110" => q_unbuf <= my_rom(3142);
      when "110001000111" => q_unbuf <= my_rom(3143);
      when "110001001000" => q_unbuf <= my_rom(3144);
      when "110001001001" => q_unbuf <= my_rom(3145);
      when "110001001010" => q_unbuf <= my_rom(3146);
      when "110001001011" => q_unbuf <= my_rom(3147);
      when "110001001100" => q_unbuf <= my_rom(3148);
      when "110001001101" => q_unbuf <= my_rom(3149);
      when "110001001110" => q_unbuf <= my_rom(3150);
      when "110001001111" => q_unbuf <= my_rom(3151);
      when "110001010000" => q_unbuf <= my_rom(3152);
      when "110001010001" => q_unbuf <= my_rom(3153);
      when "110001010010" => q_unbuf <= my_rom(3154);
      when "110001010011" => q_unbuf <= my_rom(3155);
      when "110001010100" => q_unbuf <= my_rom(3156);
      when "110001010101" => q_unbuf <= my_rom(3157);
      when "110001010110" => q_unbuf <= my_rom(3158);
      when "110001010111" => q_unbuf <= my_rom(3159);
      when "110001011000" => q_unbuf <= my_rom(3160);
      when "110001011001" => q_unbuf <= my_rom(3161);
      when "110001011010" => q_unbuf <= my_rom(3162);
      when "110001011011" => q_unbuf <= my_rom(3163);
      when "110001011100" => q_unbuf <= my_rom(3164);
      when "110001011101" => q_unbuf <= my_rom(3165);
      when "110001011110" => q_unbuf <= my_rom(3166);
      when "110001011111" => q_unbuf <= my_rom(3167);
      when "110001100000" => q_unbuf <= my_rom(3168);
      when "110001100001" => q_unbuf <= my_rom(3169);
      when "110001100010" => q_unbuf <= my_rom(3170);
      when "110001100011" => q_unbuf <= my_rom(3171);
      when "110001100100" => q_unbuf <= my_rom(3172);
      when "110001100101" => q_unbuf <= my_rom(3173);
      when "110001100110" => q_unbuf <= my_rom(3174);
      when "110001100111" => q_unbuf <= my_rom(3175);
      when "110001101000" => q_unbuf <= my_rom(3176);
      when "110001101001" => q_unbuf <= my_rom(3177);
      when "110001101010" => q_unbuf <= my_rom(3178);
      when "110001101011" => q_unbuf <= my_rom(3179);
      when "110001101100" => q_unbuf <= my_rom(3180);
      when "110001101101" => q_unbuf <= my_rom(3181);
      when "110001101110" => q_unbuf <= my_rom(3182);
      when "110001101111" => q_unbuf <= my_rom(3183);
      when "110001110000" => q_unbuf <= my_rom(3184);
      when "110001110001" => q_unbuf <= my_rom(3185);
      when "110001110010" => q_unbuf <= my_rom(3186);
      when "110001110011" => q_unbuf <= my_rom(3187);
      when "110001110100" => q_unbuf <= my_rom(3188);
      when "110001110101" => q_unbuf <= my_rom(3189);
      when "110001110110" => q_unbuf <= my_rom(3190);
      when "110001110111" => q_unbuf <= my_rom(3191);
      when "110001111000" => q_unbuf <= my_rom(3192);
      when "110001111001" => q_unbuf <= my_rom(3193);
      when "110001111010" => q_unbuf <= my_rom(3194);
      when "110001111011" => q_unbuf <= my_rom(3195);
      when "110001111100" => q_unbuf <= my_rom(3196);
      when "110001111101" => q_unbuf <= my_rom(3197);
      when "110001111110" => q_unbuf <= my_rom(3198);
      when "110001111111" => q_unbuf <= my_rom(3199);
      when "110010000000" => q_unbuf <= my_rom(3200);
      when "110010000001" => q_unbuf <= my_rom(3201);
      when "110010000010" => q_unbuf <= my_rom(3202);
      when "110010000011" => q_unbuf <= my_rom(3203);
      when "110010000100" => q_unbuf <= my_rom(3204);
      when "110010000101" => q_unbuf <= my_rom(3205);
      when "110010000110" => q_unbuf <= my_rom(3206);
      when "110010000111" => q_unbuf <= my_rom(3207);
      when "110010001000" => q_unbuf <= my_rom(3208);
      when "110010001001" => q_unbuf <= my_rom(3209);
      when "110010001010" => q_unbuf <= my_rom(3210);
      when "110010001011" => q_unbuf <= my_rom(3211);
      when "110010001100" => q_unbuf <= my_rom(3212);
      when "110010001101" => q_unbuf <= my_rom(3213);
      when "110010001110" => q_unbuf <= my_rom(3214);
      when "110010001111" => q_unbuf <= my_rom(3215);
      when "110010010000" => q_unbuf <= my_rom(3216);
      when "110010010001" => q_unbuf <= my_rom(3217);
      when "110010010010" => q_unbuf <= my_rom(3218);
      when "110010010011" => q_unbuf <= my_rom(3219);
      when "110010010100" => q_unbuf <= my_rom(3220);
      when "110010010101" => q_unbuf <= my_rom(3221);
      when "110010010110" => q_unbuf <= my_rom(3222);
      when "110010010111" => q_unbuf <= my_rom(3223);
      when "110010011000" => q_unbuf <= my_rom(3224);
      when "110010011001" => q_unbuf <= my_rom(3225);
      when "110010011010" => q_unbuf <= my_rom(3226);
      when "110010011011" => q_unbuf <= my_rom(3227);
      when "110010011100" => q_unbuf <= my_rom(3228);
      when "110010011101" => q_unbuf <= my_rom(3229);
      when "110010011110" => q_unbuf <= my_rom(3230);
      when "110010011111" => q_unbuf <= my_rom(3231);
      when "110010100000" => q_unbuf <= my_rom(3232);
      when "110010100001" => q_unbuf <= my_rom(3233);
      when "110010100010" => q_unbuf <= my_rom(3234);
      when "110010100011" => q_unbuf <= my_rom(3235);
      when "110010100100" => q_unbuf <= my_rom(3236);
      when "110010100101" => q_unbuf <= my_rom(3237);
      when "110010100110" => q_unbuf <= my_rom(3238);
      when "110010100111" => q_unbuf <= my_rom(3239);
      when "110010101000" => q_unbuf <= my_rom(3240);
      when "110010101001" => q_unbuf <= my_rom(3241);
      when "110010101010" => q_unbuf <= my_rom(3242);
      when "110010101011" => q_unbuf <= my_rom(3243);
      when "110010101100" => q_unbuf <= my_rom(3244);
      when "110010101101" => q_unbuf <= my_rom(3245);
      when "110010101110" => q_unbuf <= my_rom(3246);
      when "110010101111" => q_unbuf <= my_rom(3247);
      when "110010110000" => q_unbuf <= my_rom(3248);
      when "110010110001" => q_unbuf <= my_rom(3249);
      when "110010110010" => q_unbuf <= my_rom(3250);
      when "110010110011" => q_unbuf <= my_rom(3251);
      when "110010110100" => q_unbuf <= my_rom(3252);
      when "110010110101" => q_unbuf <= my_rom(3253);
      when "110010110110" => q_unbuf <= my_rom(3254);
      when "110010110111" => q_unbuf <= my_rom(3255);
      when "110010111000" => q_unbuf <= my_rom(3256);
      when "110010111001" => q_unbuf <= my_rom(3257);
      when "110010111010" => q_unbuf <= my_rom(3258);
      when "110010111011" => q_unbuf <= my_rom(3259);
      when "110010111100" => q_unbuf <= my_rom(3260);
      when "110010111101" => q_unbuf <= my_rom(3261);
      when "110010111110" => q_unbuf <= my_rom(3262);
      when "110010111111" => q_unbuf <= my_rom(3263);
      when "110011000000" => q_unbuf <= my_rom(3264);
      when "110011000001" => q_unbuf <= my_rom(3265);
      when "110011000010" => q_unbuf <= my_rom(3266);
      when "110011000011" => q_unbuf <= my_rom(3267);
      when "110011000100" => q_unbuf <= my_rom(3268);
      when "110011000101" => q_unbuf <= my_rom(3269);
      when "110011000110" => q_unbuf <= my_rom(3270);
      when "110011000111" => q_unbuf <= my_rom(3271);
      when "110011001000" => q_unbuf <= my_rom(3272);
      when "110011001001" => q_unbuf <= my_rom(3273);
      when "110011001010" => q_unbuf <= my_rom(3274);
      when "110011001011" => q_unbuf <= my_rom(3275);
      when "110011001100" => q_unbuf <= my_rom(3276);
      when "110011001101" => q_unbuf <= my_rom(3277);
      when "110011001110" => q_unbuf <= my_rom(3278);
      when "110011001111" => q_unbuf <= my_rom(3279);
      when "110011010000" => q_unbuf <= my_rom(3280);
      when "110011010001" => q_unbuf <= my_rom(3281);
      when "110011010010" => q_unbuf <= my_rom(3282);
      when "110011010011" => q_unbuf <= my_rom(3283);
      when "110011010100" => q_unbuf <= my_rom(3284);
      when "110011010101" => q_unbuf <= my_rom(3285);
      when "110011010110" => q_unbuf <= my_rom(3286);
      when "110011010111" => q_unbuf <= my_rom(3287);
      when "110011011000" => q_unbuf <= my_rom(3288);
      when "110011011001" => q_unbuf <= my_rom(3289);
      when "110011011010" => q_unbuf <= my_rom(3290);
      when "110011011011" => q_unbuf <= my_rom(3291);
      when "110011011100" => q_unbuf <= my_rom(3292);
      when "110011011101" => q_unbuf <= my_rom(3293);
      when "110011011110" => q_unbuf <= my_rom(3294);
      when "110011011111" => q_unbuf <= my_rom(3295);
      when "110011100000" => q_unbuf <= my_rom(3296);
      when "110011100001" => q_unbuf <= my_rom(3297);
      when "110011100010" => q_unbuf <= my_rom(3298);
      when "110011100011" => q_unbuf <= my_rom(3299);
      when "110011100100" => q_unbuf <= my_rom(3300);
      when "110011100101" => q_unbuf <= my_rom(3301);
      when "110011100110" => q_unbuf <= my_rom(3302);
      when "110011100111" => q_unbuf <= my_rom(3303);
      when "110011101000" => q_unbuf <= my_rom(3304);
      when "110011101001" => q_unbuf <= my_rom(3305);
      when "110011101010" => q_unbuf <= my_rom(3306);
      when "110011101011" => q_unbuf <= my_rom(3307);
      when "110011101100" => q_unbuf <= my_rom(3308);
      when "110011101101" => q_unbuf <= my_rom(3309);
      when "110011101110" => q_unbuf <= my_rom(3310);
      when "110011101111" => q_unbuf <= my_rom(3311);
      when "110011110000" => q_unbuf <= my_rom(3312);
      when "110011110001" => q_unbuf <= my_rom(3313);
      when "110011110010" => q_unbuf <= my_rom(3314);
      when "110011110011" => q_unbuf <= my_rom(3315);
      when "110011110100" => q_unbuf <= my_rom(3316);
      when "110011110101" => q_unbuf <= my_rom(3317);
      when "110011110110" => q_unbuf <= my_rom(3318);
      when "110011110111" => q_unbuf <= my_rom(3319);
      when "110011111000" => q_unbuf <= my_rom(3320);
      when "110011111001" => q_unbuf <= my_rom(3321);
      when "110011111010" => q_unbuf <= my_rom(3322);
      when "110011111011" => q_unbuf <= my_rom(3323);
      when "110011111100" => q_unbuf <= my_rom(3324);
      when "110011111101" => q_unbuf <= my_rom(3325);
      when "110011111110" => q_unbuf <= my_rom(3326);
      when "110011111111" => q_unbuf <= my_rom(3327);
      when "110100000000" => q_unbuf <= my_rom(3328);
      when "110100000001" => q_unbuf <= my_rom(3329);
      when "110100000010" => q_unbuf <= my_rom(3330);
      when "110100000011" => q_unbuf <= my_rom(3331);
      when "110100000100" => q_unbuf <= my_rom(3332);
      when "110100000101" => q_unbuf <= my_rom(3333);
      when "110100000110" => q_unbuf <= my_rom(3334);
      when "110100000111" => q_unbuf <= my_rom(3335);
      when "110100001000" => q_unbuf <= my_rom(3336);
      when "110100001001" => q_unbuf <= my_rom(3337);
      when "110100001010" => q_unbuf <= my_rom(3338);
      when "110100001011" => q_unbuf <= my_rom(3339);
      when "110100001100" => q_unbuf <= my_rom(3340);
      when "110100001101" => q_unbuf <= my_rom(3341);
      when "110100001110" => q_unbuf <= my_rom(3342);
      when "110100001111" => q_unbuf <= my_rom(3343);
      when "110100010000" => q_unbuf <= my_rom(3344);
      when "110100010001" => q_unbuf <= my_rom(3345);
      when "110100010010" => q_unbuf <= my_rom(3346);
      when "110100010011" => q_unbuf <= my_rom(3347);
      when "110100010100" => q_unbuf <= my_rom(3348);
      when "110100010101" => q_unbuf <= my_rom(3349);
      when "110100010110" => q_unbuf <= my_rom(3350);
      when "110100010111" => q_unbuf <= my_rom(3351);
      when "110100011000" => q_unbuf <= my_rom(3352);
      when "110100011001" => q_unbuf <= my_rom(3353);
      when "110100011010" => q_unbuf <= my_rom(3354);
      when "110100011011" => q_unbuf <= my_rom(3355);
      when "110100011100" => q_unbuf <= my_rom(3356);
      when "110100011101" => q_unbuf <= my_rom(3357);
      when "110100011110" => q_unbuf <= my_rom(3358);
      when "110100011111" => q_unbuf <= my_rom(3359);
      when "110100100000" => q_unbuf <= my_rom(3360);
      when "110100100001" => q_unbuf <= my_rom(3361);
      when "110100100010" => q_unbuf <= my_rom(3362);
      when "110100100011" => q_unbuf <= my_rom(3363);
      when "110100100100" => q_unbuf <= my_rom(3364);
      when "110100100101" => q_unbuf <= my_rom(3365);
      when "110100100110" => q_unbuf <= my_rom(3366);
      when "110100100111" => q_unbuf <= my_rom(3367);
      when "110100101000" => q_unbuf <= my_rom(3368);
      when "110100101001" => q_unbuf <= my_rom(3369);
      when "110100101010" => q_unbuf <= my_rom(3370);
      when "110100101011" => q_unbuf <= my_rom(3371);
      when "110100101100" => q_unbuf <= my_rom(3372);
      when "110100101101" => q_unbuf <= my_rom(3373);
      when "110100101110" => q_unbuf <= my_rom(3374);
      when "110100101111" => q_unbuf <= my_rom(3375);
      when "110100110000" => q_unbuf <= my_rom(3376);
      when "110100110001" => q_unbuf <= my_rom(3377);
      when "110100110010" => q_unbuf <= my_rom(3378);
      when "110100110011" => q_unbuf <= my_rom(3379);
      when "110100110100" => q_unbuf <= my_rom(3380);
      when "110100110101" => q_unbuf <= my_rom(3381);
      when "110100110110" => q_unbuf <= my_rom(3382);
      when "110100110111" => q_unbuf <= my_rom(3383);
      when "110100111000" => q_unbuf <= my_rom(3384);
      when "110100111001" => q_unbuf <= my_rom(3385);
      when "110100111010" => q_unbuf <= my_rom(3386);
      when "110100111011" => q_unbuf <= my_rom(3387);
      when "110100111100" => q_unbuf <= my_rom(3388);
      when "110100111101" => q_unbuf <= my_rom(3389);
      when "110100111110" => q_unbuf <= my_rom(3390);
      when "110100111111" => q_unbuf <= my_rom(3391);
      when "110101000000" => q_unbuf <= my_rom(3392);
      when "110101000001" => q_unbuf <= my_rom(3393);
      when "110101000010" => q_unbuf <= my_rom(3394);
      when "110101000011" => q_unbuf <= my_rom(3395);
      when "110101000100" => q_unbuf <= my_rom(3396);
      when "110101000101" => q_unbuf <= my_rom(3397);
      when "110101000110" => q_unbuf <= my_rom(3398);
      when "110101000111" => q_unbuf <= my_rom(3399);
      when "110101001000" => q_unbuf <= my_rom(3400);
      when "110101001001" => q_unbuf <= my_rom(3401);
      when "110101001010" => q_unbuf <= my_rom(3402);
      when "110101001011" => q_unbuf <= my_rom(3403);
      when "110101001100" => q_unbuf <= my_rom(3404);
      when "110101001101" => q_unbuf <= my_rom(3405);
      when "110101001110" => q_unbuf <= my_rom(3406);
      when "110101001111" => q_unbuf <= my_rom(3407);
      when "110101010000" => q_unbuf <= my_rom(3408);
      when "110101010001" => q_unbuf <= my_rom(3409);
      when "110101010010" => q_unbuf <= my_rom(3410);
      when "110101010011" => q_unbuf <= my_rom(3411);
      when "110101010100" => q_unbuf <= my_rom(3412);
      when "110101010101" => q_unbuf <= my_rom(3413);
      when "110101010110" => q_unbuf <= my_rom(3414);
      when "110101010111" => q_unbuf <= my_rom(3415);
      when "110101011000" => q_unbuf <= my_rom(3416);
      when "110101011001" => q_unbuf <= my_rom(3417);
      when "110101011010" => q_unbuf <= my_rom(3418);
      when "110101011011" => q_unbuf <= my_rom(3419);
      when "110101011100" => q_unbuf <= my_rom(3420);
      when "110101011101" => q_unbuf <= my_rom(3421);
      when "110101011110" => q_unbuf <= my_rom(3422);
      when "110101011111" => q_unbuf <= my_rom(3423);
      when "110101100000" => q_unbuf <= my_rom(3424);
      when "110101100001" => q_unbuf <= my_rom(3425);
      when "110101100010" => q_unbuf <= my_rom(3426);
      when "110101100011" => q_unbuf <= my_rom(3427);
      when "110101100100" => q_unbuf <= my_rom(3428);
      when "110101100101" => q_unbuf <= my_rom(3429);
      when "110101100110" => q_unbuf <= my_rom(3430);
      when "110101100111" => q_unbuf <= my_rom(3431);
      when "110101101000" => q_unbuf <= my_rom(3432);
      when "110101101001" => q_unbuf <= my_rom(3433);
      when "110101101010" => q_unbuf <= my_rom(3434);
      when "110101101011" => q_unbuf <= my_rom(3435);
      when "110101101100" => q_unbuf <= my_rom(3436);
      when "110101101101" => q_unbuf <= my_rom(3437);
      when "110101101110" => q_unbuf <= my_rom(3438);
      when "110101101111" => q_unbuf <= my_rom(3439);
      when "110101110000" => q_unbuf <= my_rom(3440);
      when "110101110001" => q_unbuf <= my_rom(3441);
      when "110101110010" => q_unbuf <= my_rom(3442);
      when "110101110011" => q_unbuf <= my_rom(3443);
      when "110101110100" => q_unbuf <= my_rom(3444);
      when "110101110101" => q_unbuf <= my_rom(3445);
      when "110101110110" => q_unbuf <= my_rom(3446);
      when "110101110111" => q_unbuf <= my_rom(3447);
      when "110101111000" => q_unbuf <= my_rom(3448);
      when "110101111001" => q_unbuf <= my_rom(3449);
      when "110101111010" => q_unbuf <= my_rom(3450);
      when "110101111011" => q_unbuf <= my_rom(3451);
      when "110101111100" => q_unbuf <= my_rom(3452);
      when "110101111101" => q_unbuf <= my_rom(3453);
      when "110101111110" => q_unbuf <= my_rom(3454);
      when "110101111111" => q_unbuf <= my_rom(3455);
      when "110110000000" => q_unbuf <= my_rom(3456);
      when "110110000001" => q_unbuf <= my_rom(3457);
      when "110110000010" => q_unbuf <= my_rom(3458);
      when "110110000011" => q_unbuf <= my_rom(3459);
      when "110110000100" => q_unbuf <= my_rom(3460);
      when "110110000101" => q_unbuf <= my_rom(3461);
      when "110110000110" => q_unbuf <= my_rom(3462);
      when "110110000111" => q_unbuf <= my_rom(3463);
      when "110110001000" => q_unbuf <= my_rom(3464);
      when "110110001001" => q_unbuf <= my_rom(3465);
      when "110110001010" => q_unbuf <= my_rom(3466);
      when "110110001011" => q_unbuf <= my_rom(3467);
      when "110110001100" => q_unbuf <= my_rom(3468);
      when "110110001101" => q_unbuf <= my_rom(3469);
      when "110110001110" => q_unbuf <= my_rom(3470);
      when "110110001111" => q_unbuf <= my_rom(3471);
      when "110110010000" => q_unbuf <= my_rom(3472);
      when "110110010001" => q_unbuf <= my_rom(3473);
      when "110110010010" => q_unbuf <= my_rom(3474);
      when "110110010011" => q_unbuf <= my_rom(3475);
      when "110110010100" => q_unbuf <= my_rom(3476);
      when "110110010101" => q_unbuf <= my_rom(3477);
      when "110110010110" => q_unbuf <= my_rom(3478);
      when "110110010111" => q_unbuf <= my_rom(3479);
      when "110110011000" => q_unbuf <= my_rom(3480);
      when "110110011001" => q_unbuf <= my_rom(3481);
      when "110110011010" => q_unbuf <= my_rom(3482);
      when "110110011011" => q_unbuf <= my_rom(3483);
      when "110110011100" => q_unbuf <= my_rom(3484);
      when "110110011101" => q_unbuf <= my_rom(3485);
      when "110110011110" => q_unbuf <= my_rom(3486);
      when "110110011111" => q_unbuf <= my_rom(3487);
      when "110110100000" => q_unbuf <= my_rom(3488);
      when "110110100001" => q_unbuf <= my_rom(3489);
      when "110110100010" => q_unbuf <= my_rom(3490);
      when "110110100011" => q_unbuf <= my_rom(3491);
      when "110110100100" => q_unbuf <= my_rom(3492);
      when "110110100101" => q_unbuf <= my_rom(3493);
      when "110110100110" => q_unbuf <= my_rom(3494);
      when "110110100111" => q_unbuf <= my_rom(3495);
      when "110110101000" => q_unbuf <= my_rom(3496);
      when "110110101001" => q_unbuf <= my_rom(3497);
      when "110110101010" => q_unbuf <= my_rom(3498);
      when "110110101011" => q_unbuf <= my_rom(3499);
      when "110110101100" => q_unbuf <= my_rom(3500);
      when "110110101101" => q_unbuf <= my_rom(3501);
      when "110110101110" => q_unbuf <= my_rom(3502);
      when "110110101111" => q_unbuf <= my_rom(3503);
      when "110110110000" => q_unbuf <= my_rom(3504);
      when "110110110001" => q_unbuf <= my_rom(3505);
      when "110110110010" => q_unbuf <= my_rom(3506);
      when "110110110011" => q_unbuf <= my_rom(3507);
      when "110110110100" => q_unbuf <= my_rom(3508);
      when "110110110101" => q_unbuf <= my_rom(3509);
      when "110110110110" => q_unbuf <= my_rom(3510);
      when "110110110111" => q_unbuf <= my_rom(3511);
      when "110110111000" => q_unbuf <= my_rom(3512);
      when "110110111001" => q_unbuf <= my_rom(3513);
      when "110110111010" => q_unbuf <= my_rom(3514);
      when "110110111011" => q_unbuf <= my_rom(3515);
      when "110110111100" => q_unbuf <= my_rom(3516);
      when "110110111101" => q_unbuf <= my_rom(3517);
      when "110110111110" => q_unbuf <= my_rom(3518);
      when "110110111111" => q_unbuf <= my_rom(3519);
      when "110111000000" => q_unbuf <= my_rom(3520);
      when "110111000001" => q_unbuf <= my_rom(3521);
      when "110111000010" => q_unbuf <= my_rom(3522);
      when "110111000011" => q_unbuf <= my_rom(3523);
      when "110111000100" => q_unbuf <= my_rom(3524);
      when "110111000101" => q_unbuf <= my_rom(3525);
      when "110111000110" => q_unbuf <= my_rom(3526);
      when "110111000111" => q_unbuf <= my_rom(3527);
      when "110111001000" => q_unbuf <= my_rom(3528);
      when "110111001001" => q_unbuf <= my_rom(3529);
      when "110111001010" => q_unbuf <= my_rom(3530);
      when "110111001011" => q_unbuf <= my_rom(3531);
      when "110111001100" => q_unbuf <= my_rom(3532);
      when "110111001101" => q_unbuf <= my_rom(3533);
      when "110111001110" => q_unbuf <= my_rom(3534);
      when "110111001111" => q_unbuf <= my_rom(3535);
      when "110111010000" => q_unbuf <= my_rom(3536);
      when "110111010001" => q_unbuf <= my_rom(3537);
      when "110111010010" => q_unbuf <= my_rom(3538);
      when "110111010011" => q_unbuf <= my_rom(3539);
      when "110111010100" => q_unbuf <= my_rom(3540);
      when "110111010101" => q_unbuf <= my_rom(3541);
      when "110111010110" => q_unbuf <= my_rom(3542);
      when "110111010111" => q_unbuf <= my_rom(3543);
      when "110111011000" => q_unbuf <= my_rom(3544);
      when "110111011001" => q_unbuf <= my_rom(3545);
      when "110111011010" => q_unbuf <= my_rom(3546);
      when "110111011011" => q_unbuf <= my_rom(3547);
      when "110111011100" => q_unbuf <= my_rom(3548);
      when "110111011101" => q_unbuf <= my_rom(3549);
      when "110111011110" => q_unbuf <= my_rom(3550);
      when "110111011111" => q_unbuf <= my_rom(3551);
      when "110111100000" => q_unbuf <= my_rom(3552);
      when "110111100001" => q_unbuf <= my_rom(3553);
      when "110111100010" => q_unbuf <= my_rom(3554);
      when "110111100011" => q_unbuf <= my_rom(3555);
      when "110111100100" => q_unbuf <= my_rom(3556);
      when "110111100101" => q_unbuf <= my_rom(3557);
      when "110111100110" => q_unbuf <= my_rom(3558);
      when "110111100111" => q_unbuf <= my_rom(3559);
      when "110111101000" => q_unbuf <= my_rom(3560);
      when "110111101001" => q_unbuf <= my_rom(3561);
      when "110111101010" => q_unbuf <= my_rom(3562);
      when "110111101011" => q_unbuf <= my_rom(3563);
      when "110111101100" => q_unbuf <= my_rom(3564);
      when "110111101101" => q_unbuf <= my_rom(3565);
      when "110111101110" => q_unbuf <= my_rom(3566);
      when "110111101111" => q_unbuf <= my_rom(3567);
      when "110111110000" => q_unbuf <= my_rom(3568);
      when "110111110001" => q_unbuf <= my_rom(3569);
      when "110111110010" => q_unbuf <= my_rom(3570);
      when "110111110011" => q_unbuf <= my_rom(3571);
      when "110111110100" => q_unbuf <= my_rom(3572);
      when "110111110101" => q_unbuf <= my_rom(3573);
      when "110111110110" => q_unbuf <= my_rom(3574);
      when "110111110111" => q_unbuf <= my_rom(3575);
      when "110111111000" => q_unbuf <= my_rom(3576);
      when "110111111001" => q_unbuf <= my_rom(3577);
      when "110111111010" => q_unbuf <= my_rom(3578);
      when "110111111011" => q_unbuf <= my_rom(3579);
      when "110111111100" => q_unbuf <= my_rom(3580);
      when "110111111101" => q_unbuf <= my_rom(3581);
      when "110111111110" => q_unbuf <= my_rom(3582);
      when "110111111111" => q_unbuf <= my_rom(3583);
      when "111000000000" => q_unbuf <= my_rom(3584);
      when "111000000001" => q_unbuf <= my_rom(3585);
      when "111000000010" => q_unbuf <= my_rom(3586);
      when "111000000011" => q_unbuf <= my_rom(3587);
      when "111000000100" => q_unbuf <= my_rom(3588);
      when "111000000101" => q_unbuf <= my_rom(3589);
      when "111000000110" => q_unbuf <= my_rom(3590);
      when "111000000111" => q_unbuf <= my_rom(3591);
      when "111000001000" => q_unbuf <= my_rom(3592);
      when "111000001001" => q_unbuf <= my_rom(3593);
      when "111000001010" => q_unbuf <= my_rom(3594);
      when "111000001011" => q_unbuf <= my_rom(3595);
      when "111000001100" => q_unbuf <= my_rom(3596);
      when "111000001101" => q_unbuf <= my_rom(3597);
      when "111000001110" => q_unbuf <= my_rom(3598);
      when "111000001111" => q_unbuf <= my_rom(3599);
      when "111000010000" => q_unbuf <= my_rom(3600);
      when "111000010001" => q_unbuf <= my_rom(3601);
      when "111000010010" => q_unbuf <= my_rom(3602);
      when "111000010011" => q_unbuf <= my_rom(3603);
      when "111000010100" => q_unbuf <= my_rom(3604);
      when "111000010101" => q_unbuf <= my_rom(3605);
      when "111000010110" => q_unbuf <= my_rom(3606);
      when "111000010111" => q_unbuf <= my_rom(3607);
      when "111000011000" => q_unbuf <= my_rom(3608);
      when "111000011001" => q_unbuf <= my_rom(3609);
      when "111000011010" => q_unbuf <= my_rom(3610);
      when "111000011011" => q_unbuf <= my_rom(3611);
      when "111000011100" => q_unbuf <= my_rom(3612);
      when "111000011101" => q_unbuf <= my_rom(3613);
      when "111000011110" => q_unbuf <= my_rom(3614);
      when "111000011111" => q_unbuf <= my_rom(3615);
      when "111000100000" => q_unbuf <= my_rom(3616);
      when "111000100001" => q_unbuf <= my_rom(3617);
      when "111000100010" => q_unbuf <= my_rom(3618);
      when "111000100011" => q_unbuf <= my_rom(3619);
      when "111000100100" => q_unbuf <= my_rom(3620);
      when "111000100101" => q_unbuf <= my_rom(3621);
      when "111000100110" => q_unbuf <= my_rom(3622);
      when "111000100111" => q_unbuf <= my_rom(3623);
      when "111000101000" => q_unbuf <= my_rom(3624);
      when "111000101001" => q_unbuf <= my_rom(3625);
      when "111000101010" => q_unbuf <= my_rom(3626);
      when "111000101011" => q_unbuf <= my_rom(3627);
      when "111000101100" => q_unbuf <= my_rom(3628);
      when "111000101101" => q_unbuf <= my_rom(3629);
      when "111000101110" => q_unbuf <= my_rom(3630);
      when "111000101111" => q_unbuf <= my_rom(3631);
      when "111000110000" => q_unbuf <= my_rom(3632);
      when "111000110001" => q_unbuf <= my_rom(3633);
      when "111000110010" => q_unbuf <= my_rom(3634);
      when "111000110011" => q_unbuf <= my_rom(3635);
      when "111000110100" => q_unbuf <= my_rom(3636);
      when "111000110101" => q_unbuf <= my_rom(3637);
      when "111000110110" => q_unbuf <= my_rom(3638);
      when "111000110111" => q_unbuf <= my_rom(3639);
      when "111000111000" => q_unbuf <= my_rom(3640);
      when "111000111001" => q_unbuf <= my_rom(3641);
      when "111000111010" => q_unbuf <= my_rom(3642);
      when "111000111011" => q_unbuf <= my_rom(3643);
      when "111000111100" => q_unbuf <= my_rom(3644);
      when "111000111101" => q_unbuf <= my_rom(3645);
      when "111000111110" => q_unbuf <= my_rom(3646);
      when "111000111111" => q_unbuf <= my_rom(3647);
      when "111001000000" => q_unbuf <= my_rom(3648);
      when "111001000001" => q_unbuf <= my_rom(3649);
      when "111001000010" => q_unbuf <= my_rom(3650);
      when "111001000011" => q_unbuf <= my_rom(3651);
      when "111001000100" => q_unbuf <= my_rom(3652);
      when "111001000101" => q_unbuf <= my_rom(3653);
      when "111001000110" => q_unbuf <= my_rom(3654);
      when "111001000111" => q_unbuf <= my_rom(3655);
      when "111001001000" => q_unbuf <= my_rom(3656);
      when "111001001001" => q_unbuf <= my_rom(3657);
      when "111001001010" => q_unbuf <= my_rom(3658);
      when "111001001011" => q_unbuf <= my_rom(3659);
      when "111001001100" => q_unbuf <= my_rom(3660);
      when "111001001101" => q_unbuf <= my_rom(3661);
      when "111001001110" => q_unbuf <= my_rom(3662);
      when "111001001111" => q_unbuf <= my_rom(3663);
      when "111001010000" => q_unbuf <= my_rom(3664);
      when "111001010001" => q_unbuf <= my_rom(3665);
      when "111001010010" => q_unbuf <= my_rom(3666);
      when "111001010011" => q_unbuf <= my_rom(3667);
      when "111001010100" => q_unbuf <= my_rom(3668);
      when "111001010101" => q_unbuf <= my_rom(3669);
      when "111001010110" => q_unbuf <= my_rom(3670);
      when "111001010111" => q_unbuf <= my_rom(3671);
      when "111001011000" => q_unbuf <= my_rom(3672);
      when "111001011001" => q_unbuf <= my_rom(3673);
      when "111001011010" => q_unbuf <= my_rom(3674);
      when "111001011011" => q_unbuf <= my_rom(3675);
      when "111001011100" => q_unbuf <= my_rom(3676);
      when "111001011101" => q_unbuf <= my_rom(3677);
      when "111001011110" => q_unbuf <= my_rom(3678);
      when "111001011111" => q_unbuf <= my_rom(3679);
      when "111001100000" => q_unbuf <= my_rom(3680);
      when "111001100001" => q_unbuf <= my_rom(3681);
      when "111001100010" => q_unbuf <= my_rom(3682);
      when "111001100011" => q_unbuf <= my_rom(3683);
      when "111001100100" => q_unbuf <= my_rom(3684);
      when "111001100101" => q_unbuf <= my_rom(3685);
      when "111001100110" => q_unbuf <= my_rom(3686);
      when "111001100111" => q_unbuf <= my_rom(3687);
      when "111001101000" => q_unbuf <= my_rom(3688);
      when "111001101001" => q_unbuf <= my_rom(3689);
      when "111001101010" => q_unbuf <= my_rom(3690);
      when "111001101011" => q_unbuf <= my_rom(3691);
      when "111001101100" => q_unbuf <= my_rom(3692);
      when "111001101101" => q_unbuf <= my_rom(3693);
      when "111001101110" => q_unbuf <= my_rom(3694);
      when "111001101111" => q_unbuf <= my_rom(3695);
      when "111001110000" => q_unbuf <= my_rom(3696);
      when "111001110001" => q_unbuf <= my_rom(3697);
      when "111001110010" => q_unbuf <= my_rom(3698);
      when "111001110011" => q_unbuf <= my_rom(3699);
      when "111001110100" => q_unbuf <= my_rom(3700);
      when "111001110101" => q_unbuf <= my_rom(3701);
      when "111001110110" => q_unbuf <= my_rom(3702);
      when "111001110111" => q_unbuf <= my_rom(3703);
      when "111001111000" => q_unbuf <= my_rom(3704);
      when "111001111001" => q_unbuf <= my_rom(3705);
      when "111001111010" => q_unbuf <= my_rom(3706);
      when "111001111011" => q_unbuf <= my_rom(3707);
      when "111001111100" => q_unbuf <= my_rom(3708);
      when "111001111101" => q_unbuf <= my_rom(3709);
      when "111001111110" => q_unbuf <= my_rom(3710);
      when "111001111111" => q_unbuf <= my_rom(3711);
      when "111010000000" => q_unbuf <= my_rom(3712);
      when "111010000001" => q_unbuf <= my_rom(3713);
      when "111010000010" => q_unbuf <= my_rom(3714);
      when "111010000011" => q_unbuf <= my_rom(3715);
      when "111010000100" => q_unbuf <= my_rom(3716);
      when "111010000101" => q_unbuf <= my_rom(3717);
      when "111010000110" => q_unbuf <= my_rom(3718);
      when "111010000111" => q_unbuf <= my_rom(3719);
      when "111010001000" => q_unbuf <= my_rom(3720);
      when "111010001001" => q_unbuf <= my_rom(3721);
      when "111010001010" => q_unbuf <= my_rom(3722);
      when "111010001011" => q_unbuf <= my_rom(3723);
      when "111010001100" => q_unbuf <= my_rom(3724);
      when "111010001101" => q_unbuf <= my_rom(3725);
      when "111010001110" => q_unbuf <= my_rom(3726);
      when "111010001111" => q_unbuf <= my_rom(3727);
      when "111010010000" => q_unbuf <= my_rom(3728);
      when "111010010001" => q_unbuf <= my_rom(3729);
      when "111010010010" => q_unbuf <= my_rom(3730);
      when "111010010011" => q_unbuf <= my_rom(3731);
      when "111010010100" => q_unbuf <= my_rom(3732);
      when "111010010101" => q_unbuf <= my_rom(3733);
      when "111010010110" => q_unbuf <= my_rom(3734);
      when "111010010111" => q_unbuf <= my_rom(3735);
      when "111010011000" => q_unbuf <= my_rom(3736);
      when "111010011001" => q_unbuf <= my_rom(3737);
      when "111010011010" => q_unbuf <= my_rom(3738);
      when "111010011011" => q_unbuf <= my_rom(3739);
      when "111010011100" => q_unbuf <= my_rom(3740);
      when "111010011101" => q_unbuf <= my_rom(3741);
      when "111010011110" => q_unbuf <= my_rom(3742);
      when "111010011111" => q_unbuf <= my_rom(3743);
      when "111010100000" => q_unbuf <= my_rom(3744);
      when "111010100001" => q_unbuf <= my_rom(3745);
      when "111010100010" => q_unbuf <= my_rom(3746);
      when "111010100011" => q_unbuf <= my_rom(3747);
      when "111010100100" => q_unbuf <= my_rom(3748);
      when "111010100101" => q_unbuf <= my_rom(3749);
      when "111010100110" => q_unbuf <= my_rom(3750);
      when "111010100111" => q_unbuf <= my_rom(3751);
      when "111010101000" => q_unbuf <= my_rom(3752);
      when "111010101001" => q_unbuf <= my_rom(3753);
      when "111010101010" => q_unbuf <= my_rom(3754);
      when "111010101011" => q_unbuf <= my_rom(3755);
      when "111010101100" => q_unbuf <= my_rom(3756);
      when "111010101101" => q_unbuf <= my_rom(3757);
      when "111010101110" => q_unbuf <= my_rom(3758);
      when "111010101111" => q_unbuf <= my_rom(3759);
      when "111010110000" => q_unbuf <= my_rom(3760);
      when "111010110001" => q_unbuf <= my_rom(3761);
      when "111010110010" => q_unbuf <= my_rom(3762);
      when "111010110011" => q_unbuf <= my_rom(3763);
      when "111010110100" => q_unbuf <= my_rom(3764);
      when "111010110101" => q_unbuf <= my_rom(3765);
      when "111010110110" => q_unbuf <= my_rom(3766);
      when "111010110111" => q_unbuf <= my_rom(3767);
      when "111010111000" => q_unbuf <= my_rom(3768);
      when "111010111001" => q_unbuf <= my_rom(3769);
      when "111010111010" => q_unbuf <= my_rom(3770);
      when "111010111011" => q_unbuf <= my_rom(3771);
      when "111010111100" => q_unbuf <= my_rom(3772);
      when "111010111101" => q_unbuf <= my_rom(3773);
      when "111010111110" => q_unbuf <= my_rom(3774);
      when "111010111111" => q_unbuf <= my_rom(3775);
      when "111011000000" => q_unbuf <= my_rom(3776);
      when "111011000001" => q_unbuf <= my_rom(3777);
      when "111011000010" => q_unbuf <= my_rom(3778);
      when "111011000011" => q_unbuf <= my_rom(3779);
      when "111011000100" => q_unbuf <= my_rom(3780);
      when "111011000101" => q_unbuf <= my_rom(3781);
      when "111011000110" => q_unbuf <= my_rom(3782);
      when "111011000111" => q_unbuf <= my_rom(3783);
      when "111011001000" => q_unbuf <= my_rom(3784);
      when "111011001001" => q_unbuf <= my_rom(3785);
      when "111011001010" => q_unbuf <= my_rom(3786);
      when "111011001011" => q_unbuf <= my_rom(3787);
      when "111011001100" => q_unbuf <= my_rom(3788);
      when "111011001101" => q_unbuf <= my_rom(3789);
      when "111011001110" => q_unbuf <= my_rom(3790);
      when "111011001111" => q_unbuf <= my_rom(3791);
      when "111011010000" => q_unbuf <= my_rom(3792);
      when "111011010001" => q_unbuf <= my_rom(3793);
      when "111011010010" => q_unbuf <= my_rom(3794);
      when "111011010011" => q_unbuf <= my_rom(3795);
      when "111011010100" => q_unbuf <= my_rom(3796);
      when "111011010101" => q_unbuf <= my_rom(3797);
      when "111011010110" => q_unbuf <= my_rom(3798);
      when "111011010111" => q_unbuf <= my_rom(3799);
      when "111011011000" => q_unbuf <= my_rom(3800);
      when "111011011001" => q_unbuf <= my_rom(3801);
      when "111011011010" => q_unbuf <= my_rom(3802);
      when "111011011011" => q_unbuf <= my_rom(3803);
      when "111011011100" => q_unbuf <= my_rom(3804);
      when "111011011101" => q_unbuf <= my_rom(3805);
      when "111011011110" => q_unbuf <= my_rom(3806);
      when "111011011111" => q_unbuf <= my_rom(3807);
      when "111011100000" => q_unbuf <= my_rom(3808);
      when "111011100001" => q_unbuf <= my_rom(3809);
      when "111011100010" => q_unbuf <= my_rom(3810);
      when "111011100011" => q_unbuf <= my_rom(3811);
      when "111011100100" => q_unbuf <= my_rom(3812);
      when "111011100101" => q_unbuf <= my_rom(3813);
      when "111011100110" => q_unbuf <= my_rom(3814);
      when "111011100111" => q_unbuf <= my_rom(3815);
      when "111011101000" => q_unbuf <= my_rom(3816);
      when "111011101001" => q_unbuf <= my_rom(3817);
      when "111011101010" => q_unbuf <= my_rom(3818);
      when "111011101011" => q_unbuf <= my_rom(3819);
      when "111011101100" => q_unbuf <= my_rom(3820);
      when "111011101101" => q_unbuf <= my_rom(3821);
      when "111011101110" => q_unbuf <= my_rom(3822);
      when "111011101111" => q_unbuf <= my_rom(3823);
      when "111011110000" => q_unbuf <= my_rom(3824);
      when "111011110001" => q_unbuf <= my_rom(3825);
      when "111011110010" => q_unbuf <= my_rom(3826);
      when "111011110011" => q_unbuf <= my_rom(3827);
      when "111011110100" => q_unbuf <= my_rom(3828);
      when "111011110101" => q_unbuf <= my_rom(3829);
      when "111011110110" => q_unbuf <= my_rom(3830);
      when "111011110111" => q_unbuf <= my_rom(3831);
      when "111011111000" => q_unbuf <= my_rom(3832);
      when "111011111001" => q_unbuf <= my_rom(3833);
      when "111011111010" => q_unbuf <= my_rom(3834);
      when "111011111011" => q_unbuf <= my_rom(3835);
      when "111011111100" => q_unbuf <= my_rom(3836);
      when "111011111101" => q_unbuf <= my_rom(3837);
      when "111011111110" => q_unbuf <= my_rom(3838);
      when "111011111111" => q_unbuf <= my_rom(3839);
      when "111100000000" => q_unbuf <= my_rom(3840);
      when "111100000001" => q_unbuf <= my_rom(3841);
      when "111100000010" => q_unbuf <= my_rom(3842);
      when "111100000011" => q_unbuf <= my_rom(3843);
      when "111100000100" => q_unbuf <= my_rom(3844);
      when "111100000101" => q_unbuf <= my_rom(3845);
      when "111100000110" => q_unbuf <= my_rom(3846);
      when "111100000111" => q_unbuf <= my_rom(3847);
      when "111100001000" => q_unbuf <= my_rom(3848);
      when "111100001001" => q_unbuf <= my_rom(3849);
      when "111100001010" => q_unbuf <= my_rom(3850);
      when "111100001011" => q_unbuf <= my_rom(3851);
      when "111100001100" => q_unbuf <= my_rom(3852);
      when "111100001101" => q_unbuf <= my_rom(3853);
      when "111100001110" => q_unbuf <= my_rom(3854);
      when "111100001111" => q_unbuf <= my_rom(3855);
      when "111100010000" => q_unbuf <= my_rom(3856);
      when "111100010001" => q_unbuf <= my_rom(3857);
      when "111100010010" => q_unbuf <= my_rom(3858);
      when "111100010011" => q_unbuf <= my_rom(3859);
      when "111100010100" => q_unbuf <= my_rom(3860);
      when "111100010101" => q_unbuf <= my_rom(3861);
      when "111100010110" => q_unbuf <= my_rom(3862);
      when "111100010111" => q_unbuf <= my_rom(3863);
      when "111100011000" => q_unbuf <= my_rom(3864);
      when "111100011001" => q_unbuf <= my_rom(3865);
      when "111100011010" => q_unbuf <= my_rom(3866);
      when "111100011011" => q_unbuf <= my_rom(3867);
      when "111100011100" => q_unbuf <= my_rom(3868);
      when "111100011101" => q_unbuf <= my_rom(3869);
      when "111100011110" => q_unbuf <= my_rom(3870);
      when "111100011111" => q_unbuf <= my_rom(3871);
      when "111100100000" => q_unbuf <= my_rom(3872);
      when "111100100001" => q_unbuf <= my_rom(3873);
      when "111100100010" => q_unbuf <= my_rom(3874);
      when "111100100011" => q_unbuf <= my_rom(3875);
      when "111100100100" => q_unbuf <= my_rom(3876);
      when "111100100101" => q_unbuf <= my_rom(3877);
      when "111100100110" => q_unbuf <= my_rom(3878);
      when "111100100111" => q_unbuf <= my_rom(3879);
      when "111100101000" => q_unbuf <= my_rom(3880);
      when "111100101001" => q_unbuf <= my_rom(3881);
      when "111100101010" => q_unbuf <= my_rom(3882);
      when "111100101011" => q_unbuf <= my_rom(3883);
      when "111100101100" => q_unbuf <= my_rom(3884);
      when "111100101101" => q_unbuf <= my_rom(3885);
      when "111100101110" => q_unbuf <= my_rom(3886);
      when "111100101111" => q_unbuf <= my_rom(3887);
      when "111100110000" => q_unbuf <= my_rom(3888);
      when "111100110001" => q_unbuf <= my_rom(3889);
      when "111100110010" => q_unbuf <= my_rom(3890);
      when "111100110011" => q_unbuf <= my_rom(3891);
      when "111100110100" => q_unbuf <= my_rom(3892);
      when "111100110101" => q_unbuf <= my_rom(3893);
      when "111100110110" => q_unbuf <= my_rom(3894);
      when "111100110111" => q_unbuf <= my_rom(3895);
      when "111100111000" => q_unbuf <= my_rom(3896);
      when "111100111001" => q_unbuf <= my_rom(3897);
      when "111100111010" => q_unbuf <= my_rom(3898);
      when "111100111011" => q_unbuf <= my_rom(3899);
      when "111100111100" => q_unbuf <= my_rom(3900);
      when "111100111101" => q_unbuf <= my_rom(3901);
      when "111100111110" => q_unbuf <= my_rom(3902);
      when "111100111111" => q_unbuf <= my_rom(3903);
      when "111101000000" => q_unbuf <= my_rom(3904);
      when "111101000001" => q_unbuf <= my_rom(3905);
      when "111101000010" => q_unbuf <= my_rom(3906);
      when "111101000011" => q_unbuf <= my_rom(3907);
      when "111101000100" => q_unbuf <= my_rom(3908);
      when "111101000101" => q_unbuf <= my_rom(3909);
      when "111101000110" => q_unbuf <= my_rom(3910);
      when "111101000111" => q_unbuf <= my_rom(3911);
      when "111101001000" => q_unbuf <= my_rom(3912);
      when "111101001001" => q_unbuf <= my_rom(3913);
      when "111101001010" => q_unbuf <= my_rom(3914);
      when "111101001011" => q_unbuf <= my_rom(3915);
      when "111101001100" => q_unbuf <= my_rom(3916);
      when "111101001101" => q_unbuf <= my_rom(3917);
      when "111101001110" => q_unbuf <= my_rom(3918);
      when "111101001111" => q_unbuf <= my_rom(3919);
      when "111101010000" => q_unbuf <= my_rom(3920);
      when "111101010001" => q_unbuf <= my_rom(3921);
      when "111101010010" => q_unbuf <= my_rom(3922);
      when "111101010011" => q_unbuf <= my_rom(3923);
      when "111101010100" => q_unbuf <= my_rom(3924);
      when "111101010101" => q_unbuf <= my_rom(3925);
      when "111101010110" => q_unbuf <= my_rom(3926);
      when "111101010111" => q_unbuf <= my_rom(3927);
      when "111101011000" => q_unbuf <= my_rom(3928);
      when "111101011001" => q_unbuf <= my_rom(3929);
      when "111101011010" => q_unbuf <= my_rom(3930);
      when "111101011011" => q_unbuf <= my_rom(3931);
      when "111101011100" => q_unbuf <= my_rom(3932);
      when "111101011101" => q_unbuf <= my_rom(3933);
      when "111101011110" => q_unbuf <= my_rom(3934);
      when "111101011111" => q_unbuf <= my_rom(3935);
      when "111101100000" => q_unbuf <= my_rom(3936);
      when "111101100001" => q_unbuf <= my_rom(3937);
      when "111101100010" => q_unbuf <= my_rom(3938);
      when "111101100011" => q_unbuf <= my_rom(3939);
      when "111101100100" => q_unbuf <= my_rom(3940);
      when "111101100101" => q_unbuf <= my_rom(3941);
      when "111101100110" => q_unbuf <= my_rom(3942);
      when "111101100111" => q_unbuf <= my_rom(3943);
      when "111101101000" => q_unbuf <= my_rom(3944);
      when "111101101001" => q_unbuf <= my_rom(3945);
      when "111101101010" => q_unbuf <= my_rom(3946);
      when "111101101011" => q_unbuf <= my_rom(3947);
      when "111101101100" => q_unbuf <= my_rom(3948);
      when "111101101101" => q_unbuf <= my_rom(3949);
      when "111101101110" => q_unbuf <= my_rom(3950);
      when "111101101111" => q_unbuf <= my_rom(3951);
      when "111101110000" => q_unbuf <= my_rom(3952);
      when "111101110001" => q_unbuf <= my_rom(3953);
      when "111101110010" => q_unbuf <= my_rom(3954);
      when "111101110011" => q_unbuf <= my_rom(3955);
      when "111101110100" => q_unbuf <= my_rom(3956);
      when "111101110101" => q_unbuf <= my_rom(3957);
      when "111101110110" => q_unbuf <= my_rom(3958);
      when "111101110111" => q_unbuf <= my_rom(3959);
      when "111101111000" => q_unbuf <= my_rom(3960);
      when "111101111001" => q_unbuf <= my_rom(3961);
      when "111101111010" => q_unbuf <= my_rom(3962);
      when "111101111011" => q_unbuf <= my_rom(3963);
      when "111101111100" => q_unbuf <= my_rom(3964);
      when "111101111101" => q_unbuf <= my_rom(3965);
      when "111101111110" => q_unbuf <= my_rom(3966);
      when "111101111111" => q_unbuf <= my_rom(3967);
      when "111110000000" => q_unbuf <= my_rom(3968);
      when "111110000001" => q_unbuf <= my_rom(3969);
      when "111110000010" => q_unbuf <= my_rom(3970);
      when "111110000011" => q_unbuf <= my_rom(3971);
      when "111110000100" => q_unbuf <= my_rom(3972);
      when "111110000101" => q_unbuf <= my_rom(3973);
      when "111110000110" => q_unbuf <= my_rom(3974);
      when "111110000111" => q_unbuf <= my_rom(3975);
      when "111110001000" => q_unbuf <= my_rom(3976);
      when "111110001001" => q_unbuf <= my_rom(3977);
      when "111110001010" => q_unbuf <= my_rom(3978);
      when "111110001011" => q_unbuf <= my_rom(3979);
      when "111110001100" => q_unbuf <= my_rom(3980);
      when "111110001101" => q_unbuf <= my_rom(3981);
      when "111110001110" => q_unbuf <= my_rom(3982);
      when "111110001111" => q_unbuf <= my_rom(3983);
      when "111110010000" => q_unbuf <= my_rom(3984);
      when "111110010001" => q_unbuf <= my_rom(3985);
      when "111110010010" => q_unbuf <= my_rom(3986);
      when "111110010011" => q_unbuf <= my_rom(3987);
      when "111110010100" => q_unbuf <= my_rom(3988);
      when "111110010101" => q_unbuf <= my_rom(3989);
      when "111110010110" => q_unbuf <= my_rom(3990);
      when "111110010111" => q_unbuf <= my_rom(3991);
      when "111110011000" => q_unbuf <= my_rom(3992);
      when "111110011001" => q_unbuf <= my_rom(3993);
      when "111110011010" => q_unbuf <= my_rom(3994);
      when "111110011011" => q_unbuf <= my_rom(3995);
      when "111110011100" => q_unbuf <= my_rom(3996);
      when "111110011101" => q_unbuf <= my_rom(3997);
      when "111110011110" => q_unbuf <= my_rom(3998);
      when "111110011111" => q_unbuf <= my_rom(3999);
      when "111110100000" => q_unbuf <= my_rom(4000);
      when "111110100001" => q_unbuf <= my_rom(4001);
      when "111110100010" => q_unbuf <= my_rom(4002);
      when "111110100011" => q_unbuf <= my_rom(4003);
      when "111110100100" => q_unbuf <= my_rom(4004);
      when "111110100101" => q_unbuf <= my_rom(4005);
      when "111110100110" => q_unbuf <= my_rom(4006);
      when "111110100111" => q_unbuf <= my_rom(4007);
      when "111110101000" => q_unbuf <= my_rom(4008);
      when "111110101001" => q_unbuf <= my_rom(4009);
      when "111110101010" => q_unbuf <= my_rom(4010);
      when "111110101011" => q_unbuf <= my_rom(4011);
      when "111110101100" => q_unbuf <= my_rom(4012);
      when "111110101101" => q_unbuf <= my_rom(4013);
      when "111110101110" => q_unbuf <= my_rom(4014);
      when "111110101111" => q_unbuf <= my_rom(4015);
      when "111110110000" => q_unbuf <= my_rom(4016);
      when "111110110001" => q_unbuf <= my_rom(4017);
      when "111110110010" => q_unbuf <= my_rom(4018);
      when "111110110011" => q_unbuf <= my_rom(4019);
      when "111110110100" => q_unbuf <= my_rom(4020);
      when "111110110101" => q_unbuf <= my_rom(4021);
      when "111110110110" => q_unbuf <= my_rom(4022);
      when "111110110111" => q_unbuf <= my_rom(4023);
      when "111110111000" => q_unbuf <= my_rom(4024);
      when "111110111001" => q_unbuf <= my_rom(4025);
      when "111110111010" => q_unbuf <= my_rom(4026);
      when "111110111011" => q_unbuf <= my_rom(4027);
      when "111110111100" => q_unbuf <= my_rom(4028);
      when "111110111101" => q_unbuf <= my_rom(4029);
      when "111110111110" => q_unbuf <= my_rom(4030);
      when "111110111111" => q_unbuf <= my_rom(4031);
      when "111111000000" => q_unbuf <= my_rom(4032);
      when "111111000001" => q_unbuf <= my_rom(4033);
      when "111111000010" => q_unbuf <= my_rom(4034);
      when "111111000011" => q_unbuf <= my_rom(4035);
      when "111111000100" => q_unbuf <= my_rom(4036);
      when "111111000101" => q_unbuf <= my_rom(4037);
      when "111111000110" => q_unbuf <= my_rom(4038);
      when "111111000111" => q_unbuf <= my_rom(4039);
      when "111111001000" => q_unbuf <= my_rom(4040);
      when "111111001001" => q_unbuf <= my_rom(4041);
      when "111111001010" => q_unbuf <= my_rom(4042);
      when "111111001011" => q_unbuf <= my_rom(4043);
      when "111111001100" => q_unbuf <= my_rom(4044);
      when "111111001101" => q_unbuf <= my_rom(4045);
      when "111111001110" => q_unbuf <= my_rom(4046);
      when "111111001111" => q_unbuf <= my_rom(4047);
      when "111111010000" => q_unbuf <= my_rom(4048);
      when "111111010001" => q_unbuf <= my_rom(4049);
      when "111111010010" => q_unbuf <= my_rom(4050);
      when "111111010011" => q_unbuf <= my_rom(4051);
      when "111111010100" => q_unbuf <= my_rom(4052);
      when "111111010101" => q_unbuf <= my_rom(4053);
      when "111111010110" => q_unbuf <= my_rom(4054);
      when "111111010111" => q_unbuf <= my_rom(4055);
      when "111111011000" => q_unbuf <= my_rom(4056);
      when "111111011001" => q_unbuf <= my_rom(4057);
      when "111111011010" => q_unbuf <= my_rom(4058);
      when "111111011011" => q_unbuf <= my_rom(4059);
      when "111111011100" => q_unbuf <= my_rom(4060);
      when "111111011101" => q_unbuf <= my_rom(4061);
      when "111111011110" => q_unbuf <= my_rom(4062);
      when "111111011111" => q_unbuf <= my_rom(4063);
      when "111111100000" => q_unbuf <= my_rom(4064);
      when "111111100001" => q_unbuf <= my_rom(4065);
      when "111111100010" => q_unbuf <= my_rom(4066);
      when "111111100011" => q_unbuf <= my_rom(4067);
      when "111111100100" => q_unbuf <= my_rom(4068);
      when "111111100101" => q_unbuf <= my_rom(4069);
      when "111111100110" => q_unbuf <= my_rom(4070);
      when "111111100111" => q_unbuf <= my_rom(4071);
      when "111111101000" => q_unbuf <= my_rom(4072);
      when "111111101001" => q_unbuf <= my_rom(4073);
      when "111111101010" => q_unbuf <= my_rom(4074);
      when "111111101011" => q_unbuf <= my_rom(4075);
      when "111111101100" => q_unbuf <= my_rom(4076);
      when "111111101101" => q_unbuf <= my_rom(4077);
      when "111111101110" => q_unbuf <= my_rom(4078);
      when "111111101111" => q_unbuf <= my_rom(4079);
      when "111111110000" => q_unbuf <= my_rom(4080);
      when "111111110001" => q_unbuf <= my_rom(4081);
      when "111111110010" => q_unbuf <= my_rom(4082);
      when "111111110011" => q_unbuf <= my_rom(4083);
      when "111111110100" => q_unbuf <= my_rom(4084);
      when "111111110101" => q_unbuf <= my_rom(4085);
      when "111111110110" => q_unbuf <= my_rom(4086);
      when "111111110111" => q_unbuf <= my_rom(4087);
      when "111111111000" => q_unbuf <= my_rom(4088);
      when "111111111001" => q_unbuf <= my_rom(4089);
      when "111111111010" => q_unbuf <= my_rom(4090);
      when "111111111011" => q_unbuf <= my_rom(4091);
      when "111111111100" => q_unbuf <= my_rom(4092);
      when "111111111101" => q_unbuf <= my_rom(4093);
      when "111111111110" => q_unbuf <= my_rom(4094);
      when "111111111111" => q_unbuf <= my_rom(4095);
      when others => q_unbuf <= (others => '1');
     end case;
  end process;

  process
  begin
    wait until rising_edge(clock);
    q <= q_unbuf;
  end process;

end architecture behavioral;
