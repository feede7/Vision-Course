-- Custom Vendorless ROM

library ieee;
use ieee.std_logic_1164.all;

entity lane_g_root_IP is
port (
        address : IN STD_LOGIC_VECTOR (12 DOWNTO 0);
        clock   : IN STD_LOGIC  := '1';
        q       : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
        );
end entity lane_g_root_IP;

architecture behavioral of lane_g_root_IP is
  type mem is array ( 0 to 2**13 - 1) of std_logic_vector(7 downto 0);
  constant my_Rom : mem := (
    0 => "11111111",
    1 => "11111101",
    2 => "11111011",
    3 => "11111011",
    4 => "11111010",
    5 => "11111001",
    6 => "11111001",
    7 => "11111000",
    8 => "11110111",
    9 => "11110111",
    10 => "11110111",
    11 => "11110110",
    12 => "11110110",
    13 => "11110101",
    14 => "11110101",
    15 => "11110101",
    16 => "11110100",
    17 => "11110100",
    18 => "11110011",
    19 => "11110011",
    20 => "11110011",
    21 => "11110011",
    22 => "11110010",
    23 => "11110010",
    24 => "11110010",
    25 => "11110001",
    26 => "11110001",
    27 => "11110001",
    28 => "11110001",
    29 => "11110000",
    30 => "11110000",
    31 => "11110000",
    32 => "11101111",
    33 => "11101111",
    34 => "11101111",
    35 => "11101111",
    36 => "11101111",
    37 => "11101110",
    38 => "11101110",
    39 => "11101110",
    40 => "11101110",
    41 => "11101101",
    42 => "11101101",
    43 => "11101101",
    44 => "11101101",
    45 => "11101101",
    46 => "11101100",
    47 => "11101100",
    48 => "11101100",
    49 => "11101100",
    50 => "11101011",
    51 => "11101011",
    52 => "11101011",
    53 => "11101011",
    54 => "11101011",
    55 => "11101011",
    56 => "11101010",
    57 => "11101010",
    58 => "11101010",
    59 => "11101010",
    60 => "11101010",
    61 => "11101001",
    62 => "11101001",
    63 => "11101001",
    64 => "11101001",
    65 => "11101001",
    66 => "11101001",
    67 => "11101000",
    68 => "11101000",
    69 => "11101000",
    70 => "11101000",
    71 => "11101000",
    72 => "11100111",
    73 => "11100111",
    74 => "11100111",
    75 => "11100111",
    76 => "11100111",
    77 => "11100111",
    78 => "11100111",
    79 => "11100110",
    80 => "11100110",
    81 => "11100110",
    82 => "11100110",
    83 => "11100110",
    84 => "11100110",
    85 => "11100101",
    86 => "11100101",
    87 => "11100101",
    88 => "11100101",
    89 => "11100101",
    90 => "11100101",
    91 => "11100101",
    92 => "11100100",
    93 => "11100100",
    94 => "11100100",
    95 => "11100100",
    96 => "11100100",
    97 => "11100100",
    98 => "11100011",
    99 => "11100011",
    100 => "11100011",
    101 => "11100011",
    102 => "11100011",
    103 => "11100011",
    104 => "11100011",
    105 => "11100011",
    106 => "11100010",
    107 => "11100010",
    108 => "11100010",
    109 => "11100010",
    110 => "11100010",
    111 => "11100010",
    112 => "11100010",
    113 => "11100001",
    114 => "11100001",
    115 => "11100001",
    116 => "11100001",
    117 => "11100001",
    118 => "11100001",
    119 => "11100001",
    120 => "11100001",
    121 => "11100000",
    122 => "11100000",
    123 => "11100000",
    124 => "11100000",
    125 => "11100000",
    126 => "11100000",
    127 => "11100000",
    128 => "11011111",
    129 => "11011111",
    130 => "11011111",
    131 => "11011111",
    132 => "11011111",
    133 => "11011111",
    134 => "11011111",
    135 => "11011111",
    136 => "11011111",
    137 => "11011110",
    138 => "11011110",
    139 => "11011110",
    140 => "11011110",
    141 => "11011110",
    142 => "11011110",
    143 => "11011110",
    144 => "11011110",
    145 => "11011101",
    146 => "11011101",
    147 => "11011101",
    148 => "11011101",
    149 => "11011101",
    150 => "11011101",
    151 => "11011101",
    152 => "11011101",
    153 => "11011101",
    154 => "11011100",
    155 => "11011100",
    156 => "11011100",
    157 => "11011100",
    158 => "11011100",
    159 => "11011100",
    160 => "11011100",
    161 => "11011100",
    162 => "11011011",
    163 => "11011011",
    164 => "11011011",
    165 => "11011011",
    166 => "11011011",
    167 => "11011011",
    168 => "11011011",
    169 => "11011011",
    170 => "11011011",
    171 => "11011011",
    172 => "11011010",
    173 => "11011010",
    174 => "11011010",
    175 => "11011010",
    176 => "11011010",
    177 => "11011010",
    178 => "11011010",
    179 => "11011010",
    180 => "11011010",
    181 => "11011001",
    182 => "11011001",
    183 => "11011001",
    184 => "11011001",
    185 => "11011001",
    186 => "11011001",
    187 => "11011001",
    188 => "11011001",
    189 => "11011001",
    190 => "11011001",
    191 => "11011000",
    192 => "11011000",
    193 => "11011000",
    194 => "11011000",
    195 => "11011000",
    196 => "11011000",
    197 => "11011000",
    198 => "11011000",
    199 => "11011000",
    200 => "11010111",
    201 => "11010111",
    202 => "11010111",
    203 => "11010111",
    204 => "11010111",
    205 => "11010111",
    206 => "11010111",
    207 => "11010111",
    208 => "11010111",
    209 => "11010111",
    210 => "11010111",
    211 => "11010110",
    212 => "11010110",
    213 => "11010110",
    214 => "11010110",
    215 => "11010110",
    216 => "11010110",
    217 => "11010110",
    218 => "11010110",
    219 => "11010110",
    220 => "11010110",
    221 => "11010101",
    222 => "11010101",
    223 => "11010101",
    224 => "11010101",
    225 => "11010101",
    226 => "11010101",
    227 => "11010101",
    228 => "11010101",
    229 => "11010101",
    230 => "11010101",
    231 => "11010101",
    232 => "11010100",
    233 => "11010100",
    234 => "11010100",
    235 => "11010100",
    236 => "11010100",
    237 => "11010100",
    238 => "11010100",
    239 => "11010100",
    240 => "11010100",
    241 => "11010100",
    242 => "11010011",
    243 => "11010011",
    244 => "11010011",
    245 => "11010011",
    246 => "11010011",
    247 => "11010011",
    248 => "11010011",
    249 => "11010011",
    250 => "11010011",
    251 => "11010011",
    252 => "11010011",
    253 => "11010011",
    254 => "11010010",
    255 => "11010010",
    256 => "11010010",
    257 => "11010010",
    258 => "11010010",
    259 => "11010010",
    260 => "11010010",
    261 => "11010010",
    262 => "11010010",
    263 => "11010010",
    264 => "11010010",
    265 => "11010001",
    266 => "11010001",
    267 => "11010001",
    268 => "11010001",
    269 => "11010001",
    270 => "11010001",
    271 => "11010001",
    272 => "11010001",
    273 => "11010001",
    274 => "11010001",
    275 => "11010001",
    276 => "11010001",
    277 => "11010000",
    278 => "11010000",
    279 => "11010000",
    280 => "11010000",
    281 => "11010000",
    282 => "11010000",
    283 => "11010000",
    284 => "11010000",
    285 => "11010000",
    286 => "11010000",
    287 => "11010000",
    288 => "11001111",
    289 => "11001111",
    290 => "11001111",
    291 => "11001111",
    292 => "11001111",
    293 => "11001111",
    294 => "11001111",
    295 => "11001111",
    296 => "11001111",
    297 => "11001111",
    298 => "11001111",
    299 => "11001111",
    300 => "11001111",
    301 => "11001110",
    302 => "11001110",
    303 => "11001110",
    304 => "11001110",
    305 => "11001110",
    306 => "11001110",
    307 => "11001110",
    308 => "11001110",
    309 => "11001110",
    310 => "11001110",
    311 => "11001110",
    312 => "11001110",
    313 => "11001101",
    314 => "11001101",
    315 => "11001101",
    316 => "11001101",
    317 => "11001101",
    318 => "11001101",
    319 => "11001101",
    320 => "11001101",
    321 => "11001101",
    322 => "11001101",
    323 => "11001101",
    324 => "11001101",
    325 => "11001101",
    326 => "11001100",
    327 => "11001100",
    328 => "11001100",
    329 => "11001100",
    330 => "11001100",
    331 => "11001100",
    332 => "11001100",
    333 => "11001100",
    334 => "11001100",
    335 => "11001100",
    336 => "11001100",
    337 => "11001100",
    338 => "11001011",
    339 => "11001011",
    340 => "11001011",
    341 => "11001011",
    342 => "11001011",
    343 => "11001011",
    344 => "11001011",
    345 => "11001011",
    346 => "11001011",
    347 => "11001011",
    348 => "11001011",
    349 => "11001011",
    350 => "11001011",
    351 => "11001011",
    352 => "11001010",
    353 => "11001010",
    354 => "11001010",
    355 => "11001010",
    356 => "11001010",
    357 => "11001010",
    358 => "11001010",
    359 => "11001010",
    360 => "11001010",
    361 => "11001010",
    362 => "11001010",
    363 => "11001010",
    364 => "11001010",
    365 => "11001001",
    366 => "11001001",
    367 => "11001001",
    368 => "11001001",
    369 => "11001001",
    370 => "11001001",
    371 => "11001001",
    372 => "11001001",
    373 => "11001001",
    374 => "11001001",
    375 => "11001001",
    376 => "11001001",
    377 => "11001001",
    378 => "11001001",
    379 => "11001000",
    380 => "11001000",
    381 => "11001000",
    382 => "11001000",
    383 => "11001000",
    384 => "11001000",
    385 => "11001000",
    386 => "11001000",
    387 => "11001000",
    388 => "11001000",
    389 => "11001000",
    390 => "11001000",
    391 => "11001000",
    392 => "11000111",
    393 => "11000111",
    394 => "11000111",
    395 => "11000111",
    396 => "11000111",
    397 => "11000111",
    398 => "11000111",
    399 => "11000111",
    400 => "11000111",
    401 => "11000111",
    402 => "11000111",
    403 => "11000111",
    404 => "11000111",
    405 => "11000111",
    406 => "11000111",
    407 => "11000110",
    408 => "11000110",
    409 => "11000110",
    410 => "11000110",
    411 => "11000110",
    412 => "11000110",
    413 => "11000110",
    414 => "11000110",
    415 => "11000110",
    416 => "11000110",
    417 => "11000110",
    418 => "11000110",
    419 => "11000110",
    420 => "11000110",
    421 => "11000101",
    422 => "11000101",
    423 => "11000101",
    424 => "11000101",
    425 => "11000101",
    426 => "11000101",
    427 => "11000101",
    428 => "11000101",
    429 => "11000101",
    430 => "11000101",
    431 => "11000101",
    432 => "11000101",
    433 => "11000101",
    434 => "11000101",
    435 => "11000101",
    436 => "11000100",
    437 => "11000100",
    438 => "11000100",
    439 => "11000100",
    440 => "11000100",
    441 => "11000100",
    442 => "11000100",
    443 => "11000100",
    444 => "11000100",
    445 => "11000100",
    446 => "11000100",
    447 => "11000100",
    448 => "11000100",
    449 => "11000100",
    450 => "11000011",
    451 => "11000011",
    452 => "11000011",
    453 => "11000011",
    454 => "11000011",
    455 => "11000011",
    456 => "11000011",
    457 => "11000011",
    458 => "11000011",
    459 => "11000011",
    460 => "11000011",
    461 => "11000011",
    462 => "11000011",
    463 => "11000011",
    464 => "11000011",
    465 => "11000011",
    466 => "11000010",
    467 => "11000010",
    468 => "11000010",
    469 => "11000010",
    470 => "11000010",
    471 => "11000010",
    472 => "11000010",
    473 => "11000010",
    474 => "11000010",
    475 => "11000010",
    476 => "11000010",
    477 => "11000010",
    478 => "11000010",
    479 => "11000010",
    480 => "11000010",
    481 => "11000001",
    482 => "11000001",
    483 => "11000001",
    484 => "11000001",
    485 => "11000001",
    486 => "11000001",
    487 => "11000001",
    488 => "11000001",
    489 => "11000001",
    490 => "11000001",
    491 => "11000001",
    492 => "11000001",
    493 => "11000001",
    494 => "11000001",
    495 => "11000001",
    496 => "11000001",
    497 => "11000000",
    498 => "11000000",
    499 => "11000000",
    500 => "11000000",
    501 => "11000000",
    502 => "11000000",
    503 => "11000000",
    504 => "11000000",
    505 => "11000000",
    506 => "11000000",
    507 => "11000000",
    508 => "11000000",
    509 => "11000000",
    510 => "11000000",
    511 => "11000000",
    512 => "10111111",
    513 => "10111111",
    514 => "10111111",
    515 => "10111111",
    516 => "10111111",
    517 => "10111111",
    518 => "10111111",
    519 => "10111111",
    520 => "10111111",
    521 => "10111111",
    522 => "10111111",
    523 => "10111111",
    524 => "10111111",
    525 => "10111111",
    526 => "10111111",
    527 => "10111111",
    528 => "10111111",
    529 => "10111110",
    530 => "10111110",
    531 => "10111110",
    532 => "10111110",
    533 => "10111110",
    534 => "10111110",
    535 => "10111110",
    536 => "10111110",
    537 => "10111110",
    538 => "10111110",
    539 => "10111110",
    540 => "10111110",
    541 => "10111110",
    542 => "10111110",
    543 => "10111110",
    544 => "10111110",
    545 => "10111101",
    546 => "10111101",
    547 => "10111101",
    548 => "10111101",
    549 => "10111101",
    550 => "10111101",
    551 => "10111101",
    552 => "10111101",
    553 => "10111101",
    554 => "10111101",
    555 => "10111101",
    556 => "10111101",
    557 => "10111101",
    558 => "10111101",
    559 => "10111101",
    560 => "10111101",
    561 => "10111101",
    562 => "10111100",
    563 => "10111100",
    564 => "10111100",
    565 => "10111100",
    566 => "10111100",
    567 => "10111100",
    568 => "10111100",
    569 => "10111100",
    570 => "10111100",
    571 => "10111100",
    572 => "10111100",
    573 => "10111100",
    574 => "10111100",
    575 => "10111100",
    576 => "10111100",
    577 => "10111100",
    578 => "10111011",
    579 => "10111011",
    580 => "10111011",
    581 => "10111011",
    582 => "10111011",
    583 => "10111011",
    584 => "10111011",
    585 => "10111011",
    586 => "10111011",
    587 => "10111011",
    588 => "10111011",
    589 => "10111011",
    590 => "10111011",
    591 => "10111011",
    592 => "10111011",
    593 => "10111011",
    594 => "10111011",
    595 => "10111011",
    596 => "10111010",
    597 => "10111010",
    598 => "10111010",
    599 => "10111010",
    600 => "10111010",
    601 => "10111010",
    602 => "10111010",
    603 => "10111010",
    604 => "10111010",
    605 => "10111010",
    606 => "10111010",
    607 => "10111010",
    608 => "10111010",
    609 => "10111010",
    610 => "10111010",
    611 => "10111010",
    612 => "10111010",
    613 => "10111001",
    614 => "10111001",
    615 => "10111001",
    616 => "10111001",
    617 => "10111001",
    618 => "10111001",
    619 => "10111001",
    620 => "10111001",
    621 => "10111001",
    622 => "10111001",
    623 => "10111001",
    624 => "10111001",
    625 => "10111001",
    626 => "10111001",
    627 => "10111001",
    628 => "10111001",
    629 => "10111001",
    630 => "10111001",
    631 => "10111000",
    632 => "10111000",
    633 => "10111000",
    634 => "10111000",
    635 => "10111000",
    636 => "10111000",
    637 => "10111000",
    638 => "10111000",
    639 => "10111000",
    640 => "10111000",
    641 => "10111000",
    642 => "10111000",
    643 => "10111000",
    644 => "10111000",
    645 => "10111000",
    646 => "10111000",
    647 => "10111000",
    648 => "10110111",
    649 => "10110111",
    650 => "10110111",
    651 => "10110111",
    652 => "10110111",
    653 => "10110111",
    654 => "10110111",
    655 => "10110111",
    656 => "10110111",
    657 => "10110111",
    658 => "10110111",
    659 => "10110111",
    660 => "10110111",
    661 => "10110111",
    662 => "10110111",
    663 => "10110111",
    664 => "10110111",
    665 => "10110111",
    666 => "10110111",
    667 => "10110110",
    668 => "10110110",
    669 => "10110110",
    670 => "10110110",
    671 => "10110110",
    672 => "10110110",
    673 => "10110110",
    674 => "10110110",
    675 => "10110110",
    676 => "10110110",
    677 => "10110110",
    678 => "10110110",
    679 => "10110110",
    680 => "10110110",
    681 => "10110110",
    682 => "10110110",
    683 => "10110110",
    684 => "10110110",
    685 => "10110101",
    686 => "10110101",
    687 => "10110101",
    688 => "10110101",
    689 => "10110101",
    690 => "10110101",
    691 => "10110101",
    692 => "10110101",
    693 => "10110101",
    694 => "10110101",
    695 => "10110101",
    696 => "10110101",
    697 => "10110101",
    698 => "10110101",
    699 => "10110101",
    700 => "10110101",
    701 => "10110101",
    702 => "10110101",
    703 => "10110101",
    704 => "10110100",
    705 => "10110100",
    706 => "10110100",
    707 => "10110100",
    708 => "10110100",
    709 => "10110100",
    710 => "10110100",
    711 => "10110100",
    712 => "10110100",
    713 => "10110100",
    714 => "10110100",
    715 => "10110100",
    716 => "10110100",
    717 => "10110100",
    718 => "10110100",
    719 => "10110100",
    720 => "10110100",
    721 => "10110100",
    722 => "10110011",
    723 => "10110011",
    724 => "10110011",
    725 => "10110011",
    726 => "10110011",
    727 => "10110011",
    728 => "10110011",
    729 => "10110011",
    730 => "10110011",
    731 => "10110011",
    732 => "10110011",
    733 => "10110011",
    734 => "10110011",
    735 => "10110011",
    736 => "10110011",
    737 => "10110011",
    738 => "10110011",
    739 => "10110011",
    740 => "10110011",
    741 => "10110011",
    742 => "10110010",
    743 => "10110010",
    744 => "10110010",
    745 => "10110010",
    746 => "10110010",
    747 => "10110010",
    748 => "10110010",
    749 => "10110010",
    750 => "10110010",
    751 => "10110010",
    752 => "10110010",
    753 => "10110010",
    754 => "10110010",
    755 => "10110010",
    756 => "10110010",
    757 => "10110010",
    758 => "10110010",
    759 => "10110010",
    760 => "10110010",
    761 => "10110001",
    762 => "10110001",
    763 => "10110001",
    764 => "10110001",
    765 => "10110001",
    766 => "10110001",
    767 => "10110001",
    768 => "10110001",
    769 => "10110001",
    770 => "10110001",
    771 => "10110001",
    772 => "10110001",
    773 => "10110001",
    774 => "10110001",
    775 => "10110001",
    776 => "10110001",
    777 => "10110001",
    778 => "10110001",
    779 => "10110001",
    780 => "10110001",
    781 => "10110000",
    782 => "10110000",
    783 => "10110000",
    784 => "10110000",
    785 => "10110000",
    786 => "10110000",
    787 => "10110000",
    788 => "10110000",
    789 => "10110000",
    790 => "10110000",
    791 => "10110000",
    792 => "10110000",
    793 => "10110000",
    794 => "10110000",
    795 => "10110000",
    796 => "10110000",
    797 => "10110000",
    798 => "10110000",
    799 => "10110000",
    800 => "10101111",
    801 => "10101111",
    802 => "10101111",
    803 => "10101111",
    804 => "10101111",
    805 => "10101111",
    806 => "10101111",
    807 => "10101111",
    808 => "10101111",
    809 => "10101111",
    810 => "10101111",
    811 => "10101111",
    812 => "10101111",
    813 => "10101111",
    814 => "10101111",
    815 => "10101111",
    816 => "10101111",
    817 => "10101111",
    818 => "10101111",
    819 => "10101111",
    820 => "10101111",
    821 => "10101110",
    822 => "10101110",
    823 => "10101110",
    824 => "10101110",
    825 => "10101110",
    826 => "10101110",
    827 => "10101110",
    828 => "10101110",
    829 => "10101110",
    830 => "10101110",
    831 => "10101110",
    832 => "10101110",
    833 => "10101110",
    834 => "10101110",
    835 => "10101110",
    836 => "10101110",
    837 => "10101110",
    838 => "10101110",
    839 => "10101110",
    840 => "10101110",
    841 => "10101101",
    842 => "10101101",
    843 => "10101101",
    844 => "10101101",
    845 => "10101101",
    846 => "10101101",
    847 => "10101101",
    848 => "10101101",
    849 => "10101101",
    850 => "10101101",
    851 => "10101101",
    852 => "10101101",
    853 => "10101101",
    854 => "10101101",
    855 => "10101101",
    856 => "10101101",
    857 => "10101101",
    858 => "10101101",
    859 => "10101101",
    860 => "10101101",
    861 => "10101101",
    862 => "10101100",
    863 => "10101100",
    864 => "10101100",
    865 => "10101100",
    866 => "10101100",
    867 => "10101100",
    868 => "10101100",
    869 => "10101100",
    870 => "10101100",
    871 => "10101100",
    872 => "10101100",
    873 => "10101100",
    874 => "10101100",
    875 => "10101100",
    876 => "10101100",
    877 => "10101100",
    878 => "10101100",
    879 => "10101100",
    880 => "10101100",
    881 => "10101100",
    882 => "10101011",
    883 => "10101011",
    884 => "10101011",
    885 => "10101011",
    886 => "10101011",
    887 => "10101011",
    888 => "10101011",
    889 => "10101011",
    890 => "10101011",
    891 => "10101011",
    892 => "10101011",
    893 => "10101011",
    894 => "10101011",
    895 => "10101011",
    896 => "10101011",
    897 => "10101011",
    898 => "10101011",
    899 => "10101011",
    900 => "10101011",
    901 => "10101011",
    902 => "10101011",
    903 => "10101011",
    904 => "10101010",
    905 => "10101010",
    906 => "10101010",
    907 => "10101010",
    908 => "10101010",
    909 => "10101010",
    910 => "10101010",
    911 => "10101010",
    912 => "10101010",
    913 => "10101010",
    914 => "10101010",
    915 => "10101010",
    916 => "10101010",
    917 => "10101010",
    918 => "10101010",
    919 => "10101010",
    920 => "10101010",
    921 => "10101010",
    922 => "10101010",
    923 => "10101010",
    924 => "10101010",
    925 => "10101001",
    926 => "10101001",
    927 => "10101001",
    928 => "10101001",
    929 => "10101001",
    930 => "10101001",
    931 => "10101001",
    932 => "10101001",
    933 => "10101001",
    934 => "10101001",
    935 => "10101001",
    936 => "10101001",
    937 => "10101001",
    938 => "10101001",
    939 => "10101001",
    940 => "10101001",
    941 => "10101001",
    942 => "10101001",
    943 => "10101001",
    944 => "10101001",
    945 => "10101001",
    946 => "10101001",
    947 => "10101000",
    948 => "10101000",
    949 => "10101000",
    950 => "10101000",
    951 => "10101000",
    952 => "10101000",
    953 => "10101000",
    954 => "10101000",
    955 => "10101000",
    956 => "10101000",
    957 => "10101000",
    958 => "10101000",
    959 => "10101000",
    960 => "10101000",
    961 => "10101000",
    962 => "10101000",
    963 => "10101000",
    964 => "10101000",
    965 => "10101000",
    966 => "10101000",
    967 => "10101000",
    968 => "10100111",
    969 => "10100111",
    970 => "10100111",
    971 => "10100111",
    972 => "10100111",
    973 => "10100111",
    974 => "10100111",
    975 => "10100111",
    976 => "10100111",
    977 => "10100111",
    978 => "10100111",
    979 => "10100111",
    980 => "10100111",
    981 => "10100111",
    982 => "10100111",
    983 => "10100111",
    984 => "10100111",
    985 => "10100111",
    986 => "10100111",
    987 => "10100111",
    988 => "10100111",
    989 => "10100111",
    990 => "10100111",
    991 => "10100110",
    992 => "10100110",
    993 => "10100110",
    994 => "10100110",
    995 => "10100110",
    996 => "10100110",
    997 => "10100110",
    998 => "10100110",
    999 => "10100110",
    1000 => "10100110",
    1001 => "10100110",
    1002 => "10100110",
    1003 => "10100110",
    1004 => "10100110",
    1005 => "10100110",
    1006 => "10100110",
    1007 => "10100110",
    1008 => "10100110",
    1009 => "10100110",
    1010 => "10100110",
    1011 => "10100110",
    1012 => "10100110",
    1013 => "10100101",
    1014 => "10100101",
    1015 => "10100101",
    1016 => "10100101",
    1017 => "10100101",
    1018 => "10100101",
    1019 => "10100101",
    1020 => "10100101",
    1021 => "10100101",
    1022 => "10100101",
    1023 => "10100101",
    1024 => "10100101",
    1025 => "10100101",
    1026 => "10100101",
    1027 => "10100101",
    1028 => "10100101",
    1029 => "10100101",
    1030 => "10100101",
    1031 => "10100101",
    1032 => "10100101",
    1033 => "10100101",
    1034 => "10100101",
    1035 => "10100101",
    1036 => "10100100",
    1037 => "10100100",
    1038 => "10100100",
    1039 => "10100100",
    1040 => "10100100",
    1041 => "10100100",
    1042 => "10100100",
    1043 => "10100100",
    1044 => "10100100",
    1045 => "10100100",
    1046 => "10100100",
    1047 => "10100100",
    1048 => "10100100",
    1049 => "10100100",
    1050 => "10100100",
    1051 => "10100100",
    1052 => "10100100",
    1053 => "10100100",
    1054 => "10100100",
    1055 => "10100100",
    1056 => "10100100",
    1057 => "10100100",
    1058 => "10100011",
    1059 => "10100011",
    1060 => "10100011",
    1061 => "10100011",
    1062 => "10100011",
    1063 => "10100011",
    1064 => "10100011",
    1065 => "10100011",
    1066 => "10100011",
    1067 => "10100011",
    1068 => "10100011",
    1069 => "10100011",
    1070 => "10100011",
    1071 => "10100011",
    1072 => "10100011",
    1073 => "10100011",
    1074 => "10100011",
    1075 => "10100011",
    1076 => "10100011",
    1077 => "10100011",
    1078 => "10100011",
    1079 => "10100011",
    1080 => "10100011",
    1081 => "10100011",
    1082 => "10100010",
    1083 => "10100010",
    1084 => "10100010",
    1085 => "10100010",
    1086 => "10100010",
    1087 => "10100010",
    1088 => "10100010",
    1089 => "10100010",
    1090 => "10100010",
    1091 => "10100010",
    1092 => "10100010",
    1093 => "10100010",
    1094 => "10100010",
    1095 => "10100010",
    1096 => "10100010",
    1097 => "10100010",
    1098 => "10100010",
    1099 => "10100010",
    1100 => "10100010",
    1101 => "10100010",
    1102 => "10100010",
    1103 => "10100010",
    1104 => "10100010",
    1105 => "10100001",
    1106 => "10100001",
    1107 => "10100001",
    1108 => "10100001",
    1109 => "10100001",
    1110 => "10100001",
    1111 => "10100001",
    1112 => "10100001",
    1113 => "10100001",
    1114 => "10100001",
    1115 => "10100001",
    1116 => "10100001",
    1117 => "10100001",
    1118 => "10100001",
    1119 => "10100001",
    1120 => "10100001",
    1121 => "10100001",
    1122 => "10100001",
    1123 => "10100001",
    1124 => "10100001",
    1125 => "10100001",
    1126 => "10100001",
    1127 => "10100001",
    1128 => "10100001",
    1129 => "10100000",
    1130 => "10100000",
    1131 => "10100000",
    1132 => "10100000",
    1133 => "10100000",
    1134 => "10100000",
    1135 => "10100000",
    1136 => "10100000",
    1137 => "10100000",
    1138 => "10100000",
    1139 => "10100000",
    1140 => "10100000",
    1141 => "10100000",
    1142 => "10100000",
    1143 => "10100000",
    1144 => "10100000",
    1145 => "10100000",
    1146 => "10100000",
    1147 => "10100000",
    1148 => "10100000",
    1149 => "10100000",
    1150 => "10100000",
    1151 => "10100000",
    1152 => "10011111",
    1153 => "10011111",
    1154 => "10011111",
    1155 => "10011111",
    1156 => "10011111",
    1157 => "10011111",
    1158 => "10011111",
    1159 => "10011111",
    1160 => "10011111",
    1161 => "10011111",
    1162 => "10011111",
    1163 => "10011111",
    1164 => "10011111",
    1165 => "10011111",
    1166 => "10011111",
    1167 => "10011111",
    1168 => "10011111",
    1169 => "10011111",
    1170 => "10011111",
    1171 => "10011111",
    1172 => "10011111",
    1173 => "10011111",
    1174 => "10011111",
    1175 => "10011111",
    1176 => "10011111",
    1177 => "10011110",
    1178 => "10011110",
    1179 => "10011110",
    1180 => "10011110",
    1181 => "10011110",
    1182 => "10011110",
    1183 => "10011110",
    1184 => "10011110",
    1185 => "10011110",
    1186 => "10011110",
    1187 => "10011110",
    1188 => "10011110",
    1189 => "10011110",
    1190 => "10011110",
    1191 => "10011110",
    1192 => "10011110",
    1193 => "10011110",
    1194 => "10011110",
    1195 => "10011110",
    1196 => "10011110",
    1197 => "10011110",
    1198 => "10011110",
    1199 => "10011110",
    1200 => "10011110",
    1201 => "10011101",
    1202 => "10011101",
    1203 => "10011101",
    1204 => "10011101",
    1205 => "10011101",
    1206 => "10011101",
    1207 => "10011101",
    1208 => "10011101",
    1209 => "10011101",
    1210 => "10011101",
    1211 => "10011101",
    1212 => "10011101",
    1213 => "10011101",
    1214 => "10011101",
    1215 => "10011101",
    1216 => "10011101",
    1217 => "10011101",
    1218 => "10011101",
    1219 => "10011101",
    1220 => "10011101",
    1221 => "10011101",
    1222 => "10011101",
    1223 => "10011101",
    1224 => "10011101",
    1225 => "10011101",
    1226 => "10011100",
    1227 => "10011100",
    1228 => "10011100",
    1229 => "10011100",
    1230 => "10011100",
    1231 => "10011100",
    1232 => "10011100",
    1233 => "10011100",
    1234 => "10011100",
    1235 => "10011100",
    1236 => "10011100",
    1237 => "10011100",
    1238 => "10011100",
    1239 => "10011100",
    1240 => "10011100",
    1241 => "10011100",
    1242 => "10011100",
    1243 => "10011100",
    1244 => "10011100",
    1245 => "10011100",
    1246 => "10011100",
    1247 => "10011100",
    1248 => "10011100",
    1249 => "10011100",
    1250 => "10011011",
    1251 => "10011011",
    1252 => "10011011",
    1253 => "10011011",
    1254 => "10011011",
    1255 => "10011011",
    1256 => "10011011",
    1257 => "10011011",
    1258 => "10011011",
    1259 => "10011011",
    1260 => "10011011",
    1261 => "10011011",
    1262 => "10011011",
    1263 => "10011011",
    1264 => "10011011",
    1265 => "10011011",
    1266 => "10011011",
    1267 => "10011011",
    1268 => "10011011",
    1269 => "10011011",
    1270 => "10011011",
    1271 => "10011011",
    1272 => "10011011",
    1273 => "10011011",
    1274 => "10011011",
    1275 => "10011011",
    1276 => "10011010",
    1277 => "10011010",
    1278 => "10011010",
    1279 => "10011010",
    1280 => "10011010",
    1281 => "10011010",
    1282 => "10011010",
    1283 => "10011010",
    1284 => "10011010",
    1285 => "10011010",
    1286 => "10011010",
    1287 => "10011010",
    1288 => "10011010",
    1289 => "10011010",
    1290 => "10011010",
    1291 => "10011010",
    1292 => "10011010",
    1293 => "10011010",
    1294 => "10011010",
    1295 => "10011010",
    1296 => "10011010",
    1297 => "10011010",
    1298 => "10011010",
    1299 => "10011010",
    1300 => "10011010",
    1301 => "10011001",
    1302 => "10011001",
    1303 => "10011001",
    1304 => "10011001",
    1305 => "10011001",
    1306 => "10011001",
    1307 => "10011001",
    1308 => "10011001",
    1309 => "10011001",
    1310 => "10011001",
    1311 => "10011001",
    1312 => "10011001",
    1313 => "10011001",
    1314 => "10011001",
    1315 => "10011001",
    1316 => "10011001",
    1317 => "10011001",
    1318 => "10011001",
    1319 => "10011001",
    1320 => "10011001",
    1321 => "10011001",
    1322 => "10011001",
    1323 => "10011001",
    1324 => "10011001",
    1325 => "10011001",
    1326 => "10011001",
    1327 => "10011000",
    1328 => "10011000",
    1329 => "10011000",
    1330 => "10011000",
    1331 => "10011000",
    1332 => "10011000",
    1333 => "10011000",
    1334 => "10011000",
    1335 => "10011000",
    1336 => "10011000",
    1337 => "10011000",
    1338 => "10011000",
    1339 => "10011000",
    1340 => "10011000",
    1341 => "10011000",
    1342 => "10011000",
    1343 => "10011000",
    1344 => "10011000",
    1345 => "10011000",
    1346 => "10011000",
    1347 => "10011000",
    1348 => "10011000",
    1349 => "10011000",
    1350 => "10011000",
    1351 => "10011000",
    1352 => "10010111",
    1353 => "10010111",
    1354 => "10010111",
    1355 => "10010111",
    1356 => "10010111",
    1357 => "10010111",
    1358 => "10010111",
    1359 => "10010111",
    1360 => "10010111",
    1361 => "10010111",
    1362 => "10010111",
    1363 => "10010111",
    1364 => "10010111",
    1365 => "10010111",
    1366 => "10010111",
    1367 => "10010111",
    1368 => "10010111",
    1369 => "10010111",
    1370 => "10010111",
    1371 => "10010111",
    1372 => "10010111",
    1373 => "10010111",
    1374 => "10010111",
    1375 => "10010111",
    1376 => "10010111",
    1377 => "10010111",
    1378 => "10010111",
    1379 => "10010110",
    1380 => "10010110",
    1381 => "10010110",
    1382 => "10010110",
    1383 => "10010110",
    1384 => "10010110",
    1385 => "10010110",
    1386 => "10010110",
    1387 => "10010110",
    1388 => "10010110",
    1389 => "10010110",
    1390 => "10010110",
    1391 => "10010110",
    1392 => "10010110",
    1393 => "10010110",
    1394 => "10010110",
    1395 => "10010110",
    1396 => "10010110",
    1397 => "10010110",
    1398 => "10010110",
    1399 => "10010110",
    1400 => "10010110",
    1401 => "10010110",
    1402 => "10010110",
    1403 => "10010110",
    1404 => "10010110",
    1405 => "10010101",
    1406 => "10010101",
    1407 => "10010101",
    1408 => "10010101",
    1409 => "10010101",
    1410 => "10010101",
    1411 => "10010101",
    1412 => "10010101",
    1413 => "10010101",
    1414 => "10010101",
    1415 => "10010101",
    1416 => "10010101",
    1417 => "10010101",
    1418 => "10010101",
    1419 => "10010101",
    1420 => "10010101",
    1421 => "10010101",
    1422 => "10010101",
    1423 => "10010101",
    1424 => "10010101",
    1425 => "10010101",
    1426 => "10010101",
    1427 => "10010101",
    1428 => "10010101",
    1429 => "10010101",
    1430 => "10010101",
    1431 => "10010101",
    1432 => "10010100",
    1433 => "10010100",
    1434 => "10010100",
    1435 => "10010100",
    1436 => "10010100",
    1437 => "10010100",
    1438 => "10010100",
    1439 => "10010100",
    1440 => "10010100",
    1441 => "10010100",
    1442 => "10010100",
    1443 => "10010100",
    1444 => "10010100",
    1445 => "10010100",
    1446 => "10010100",
    1447 => "10010100",
    1448 => "10010100",
    1449 => "10010100",
    1450 => "10010100",
    1451 => "10010100",
    1452 => "10010100",
    1453 => "10010100",
    1454 => "10010100",
    1455 => "10010100",
    1456 => "10010100",
    1457 => "10010100",
    1458 => "10010011",
    1459 => "10010011",
    1460 => "10010011",
    1461 => "10010011",
    1462 => "10010011",
    1463 => "10010011",
    1464 => "10010011",
    1465 => "10010011",
    1466 => "10010011",
    1467 => "10010011",
    1468 => "10010011",
    1469 => "10010011",
    1470 => "10010011",
    1471 => "10010011",
    1472 => "10010011",
    1473 => "10010011",
    1474 => "10010011",
    1475 => "10010011",
    1476 => "10010011",
    1477 => "10010011",
    1478 => "10010011",
    1479 => "10010011",
    1480 => "10010011",
    1481 => "10010011",
    1482 => "10010011",
    1483 => "10010011",
    1484 => "10010011",
    1485 => "10010011",
    1486 => "10010010",
    1487 => "10010010",
    1488 => "10010010",
    1489 => "10010010",
    1490 => "10010010",
    1491 => "10010010",
    1492 => "10010010",
    1493 => "10010010",
    1494 => "10010010",
    1495 => "10010010",
    1496 => "10010010",
    1497 => "10010010",
    1498 => "10010010",
    1499 => "10010010",
    1500 => "10010010",
    1501 => "10010010",
    1502 => "10010010",
    1503 => "10010010",
    1504 => "10010010",
    1505 => "10010010",
    1506 => "10010010",
    1507 => "10010010",
    1508 => "10010010",
    1509 => "10010010",
    1510 => "10010010",
    1511 => "10010010",
    1512 => "10010010",
    1513 => "10010001",
    1514 => "10010001",
    1515 => "10010001",
    1516 => "10010001",
    1517 => "10010001",
    1518 => "10010001",
    1519 => "10010001",
    1520 => "10010001",
    1521 => "10010001",
    1522 => "10010001",
    1523 => "10010001",
    1524 => "10010001",
    1525 => "10010001",
    1526 => "10010001",
    1527 => "10010001",
    1528 => "10010001",
    1529 => "10010001",
    1530 => "10010001",
    1531 => "10010001",
    1532 => "10010001",
    1533 => "10010001",
    1534 => "10010001",
    1535 => "10010001",
    1536 => "10010001",
    1537 => "10010001",
    1538 => "10010001",
    1539 => "10010001",
    1540 => "10010001",
    1541 => "10010000",
    1542 => "10010000",
    1543 => "10010000",
    1544 => "10010000",
    1545 => "10010000",
    1546 => "10010000",
    1547 => "10010000",
    1548 => "10010000",
    1549 => "10010000",
    1550 => "10010000",
    1551 => "10010000",
    1552 => "10010000",
    1553 => "10010000",
    1554 => "10010000",
    1555 => "10010000",
    1556 => "10010000",
    1557 => "10010000",
    1558 => "10010000",
    1559 => "10010000",
    1560 => "10010000",
    1561 => "10010000",
    1562 => "10010000",
    1563 => "10010000",
    1564 => "10010000",
    1565 => "10010000",
    1566 => "10010000",
    1567 => "10010000",
    1568 => "10001111",
    1569 => "10001111",
    1570 => "10001111",
    1571 => "10001111",
    1572 => "10001111",
    1573 => "10001111",
    1574 => "10001111",
    1575 => "10001111",
    1576 => "10001111",
    1577 => "10001111",
    1578 => "10001111",
    1579 => "10001111",
    1580 => "10001111",
    1581 => "10001111",
    1582 => "10001111",
    1583 => "10001111",
    1584 => "10001111",
    1585 => "10001111",
    1586 => "10001111",
    1587 => "10001111",
    1588 => "10001111",
    1589 => "10001111",
    1590 => "10001111",
    1591 => "10001111",
    1592 => "10001111",
    1593 => "10001111",
    1594 => "10001111",
    1595 => "10001111",
    1596 => "10001111",
    1597 => "10001110",
    1598 => "10001110",
    1599 => "10001110",
    1600 => "10001110",
    1601 => "10001110",
    1602 => "10001110",
    1603 => "10001110",
    1604 => "10001110",
    1605 => "10001110",
    1606 => "10001110",
    1607 => "10001110",
    1608 => "10001110",
    1609 => "10001110",
    1610 => "10001110",
    1611 => "10001110",
    1612 => "10001110",
    1613 => "10001110",
    1614 => "10001110",
    1615 => "10001110",
    1616 => "10001110",
    1617 => "10001110",
    1618 => "10001110",
    1619 => "10001110",
    1620 => "10001110",
    1621 => "10001110",
    1622 => "10001110",
    1623 => "10001110",
    1624 => "10001110",
    1625 => "10001101",
    1626 => "10001101",
    1627 => "10001101",
    1628 => "10001101",
    1629 => "10001101",
    1630 => "10001101",
    1631 => "10001101",
    1632 => "10001101",
    1633 => "10001101",
    1634 => "10001101",
    1635 => "10001101",
    1636 => "10001101",
    1637 => "10001101",
    1638 => "10001101",
    1639 => "10001101",
    1640 => "10001101",
    1641 => "10001101",
    1642 => "10001101",
    1643 => "10001101",
    1644 => "10001101",
    1645 => "10001101",
    1646 => "10001101",
    1647 => "10001101",
    1648 => "10001101",
    1649 => "10001101",
    1650 => "10001101",
    1651 => "10001101",
    1652 => "10001101",
    1653 => "10001101",
    1654 => "10001100",
    1655 => "10001100",
    1656 => "10001100",
    1657 => "10001100",
    1658 => "10001100",
    1659 => "10001100",
    1660 => "10001100",
    1661 => "10001100",
    1662 => "10001100",
    1663 => "10001100",
    1664 => "10001100",
    1665 => "10001100",
    1666 => "10001100",
    1667 => "10001100",
    1668 => "10001100",
    1669 => "10001100",
    1670 => "10001100",
    1671 => "10001100",
    1672 => "10001100",
    1673 => "10001100",
    1674 => "10001100",
    1675 => "10001100",
    1676 => "10001100",
    1677 => "10001100",
    1678 => "10001100",
    1679 => "10001100",
    1680 => "10001100",
    1681 => "10001100",
    1682 => "10001011",
    1683 => "10001011",
    1684 => "10001011",
    1685 => "10001011",
    1686 => "10001011",
    1687 => "10001011",
    1688 => "10001011",
    1689 => "10001011",
    1690 => "10001011",
    1691 => "10001011",
    1692 => "10001011",
    1693 => "10001011",
    1694 => "10001011",
    1695 => "10001011",
    1696 => "10001011",
    1697 => "10001011",
    1698 => "10001011",
    1699 => "10001011",
    1700 => "10001011",
    1701 => "10001011",
    1702 => "10001011",
    1703 => "10001011",
    1704 => "10001011",
    1705 => "10001011",
    1706 => "10001011",
    1707 => "10001011",
    1708 => "10001011",
    1709 => "10001011",
    1710 => "10001011",
    1711 => "10001011",
    1712 => "10001010",
    1713 => "10001010",
    1714 => "10001010",
    1715 => "10001010",
    1716 => "10001010",
    1717 => "10001010",
    1718 => "10001010",
    1719 => "10001010",
    1720 => "10001010",
    1721 => "10001010",
    1722 => "10001010",
    1723 => "10001010",
    1724 => "10001010",
    1725 => "10001010",
    1726 => "10001010",
    1727 => "10001010",
    1728 => "10001010",
    1729 => "10001010",
    1730 => "10001010",
    1731 => "10001010",
    1732 => "10001010",
    1733 => "10001010",
    1734 => "10001010",
    1735 => "10001010",
    1736 => "10001010",
    1737 => "10001010",
    1738 => "10001010",
    1739 => "10001010",
    1740 => "10001010",
    1741 => "10001001",
    1742 => "10001001",
    1743 => "10001001",
    1744 => "10001001",
    1745 => "10001001",
    1746 => "10001001",
    1747 => "10001001",
    1748 => "10001001",
    1749 => "10001001",
    1750 => "10001001",
    1751 => "10001001",
    1752 => "10001001",
    1753 => "10001001",
    1754 => "10001001",
    1755 => "10001001",
    1756 => "10001001",
    1757 => "10001001",
    1758 => "10001001",
    1759 => "10001001",
    1760 => "10001001",
    1761 => "10001001",
    1762 => "10001001",
    1763 => "10001001",
    1764 => "10001001",
    1765 => "10001001",
    1766 => "10001001",
    1767 => "10001001",
    1768 => "10001001",
    1769 => "10001001",
    1770 => "10001001",
    1771 => "10001000",
    1772 => "10001000",
    1773 => "10001000",
    1774 => "10001000",
    1775 => "10001000",
    1776 => "10001000",
    1777 => "10001000",
    1778 => "10001000",
    1779 => "10001000",
    1780 => "10001000",
    1781 => "10001000",
    1782 => "10001000",
    1783 => "10001000",
    1784 => "10001000",
    1785 => "10001000",
    1786 => "10001000",
    1787 => "10001000",
    1788 => "10001000",
    1789 => "10001000",
    1790 => "10001000",
    1791 => "10001000",
    1792 => "10001000",
    1793 => "10001000",
    1794 => "10001000",
    1795 => "10001000",
    1796 => "10001000",
    1797 => "10001000",
    1798 => "10001000",
    1799 => "10001000",
    1800 => "10000111",
    1801 => "10000111",
    1802 => "10000111",
    1803 => "10000111",
    1804 => "10000111",
    1805 => "10000111",
    1806 => "10000111",
    1807 => "10000111",
    1808 => "10000111",
    1809 => "10000111",
    1810 => "10000111",
    1811 => "10000111",
    1812 => "10000111",
    1813 => "10000111",
    1814 => "10000111",
    1815 => "10000111",
    1816 => "10000111",
    1817 => "10000111",
    1818 => "10000111",
    1819 => "10000111",
    1820 => "10000111",
    1821 => "10000111",
    1822 => "10000111",
    1823 => "10000111",
    1824 => "10000111",
    1825 => "10000111",
    1826 => "10000111",
    1827 => "10000111",
    1828 => "10000111",
    1829 => "10000111",
    1830 => "10000111",
    1831 => "10000110",
    1832 => "10000110",
    1833 => "10000110",
    1834 => "10000110",
    1835 => "10000110",
    1836 => "10000110",
    1837 => "10000110",
    1838 => "10000110",
    1839 => "10000110",
    1840 => "10000110",
    1841 => "10000110",
    1842 => "10000110",
    1843 => "10000110",
    1844 => "10000110",
    1845 => "10000110",
    1846 => "10000110",
    1847 => "10000110",
    1848 => "10000110",
    1849 => "10000110",
    1850 => "10000110",
    1851 => "10000110",
    1852 => "10000110",
    1853 => "10000110",
    1854 => "10000110",
    1855 => "10000110",
    1856 => "10000110",
    1857 => "10000110",
    1858 => "10000110",
    1859 => "10000110",
    1860 => "10000110",
    1861 => "10000101",
    1862 => "10000101",
    1863 => "10000101",
    1864 => "10000101",
    1865 => "10000101",
    1866 => "10000101",
    1867 => "10000101",
    1868 => "10000101",
    1869 => "10000101",
    1870 => "10000101",
    1871 => "10000101",
    1872 => "10000101",
    1873 => "10000101",
    1874 => "10000101",
    1875 => "10000101",
    1876 => "10000101",
    1877 => "10000101",
    1878 => "10000101",
    1879 => "10000101",
    1880 => "10000101",
    1881 => "10000101",
    1882 => "10000101",
    1883 => "10000101",
    1884 => "10000101",
    1885 => "10000101",
    1886 => "10000101",
    1887 => "10000101",
    1888 => "10000101",
    1889 => "10000101",
    1890 => "10000101",
    1891 => "10000101",
    1892 => "10000100",
    1893 => "10000100",
    1894 => "10000100",
    1895 => "10000100",
    1896 => "10000100",
    1897 => "10000100",
    1898 => "10000100",
    1899 => "10000100",
    1900 => "10000100",
    1901 => "10000100",
    1902 => "10000100",
    1903 => "10000100",
    1904 => "10000100",
    1905 => "10000100",
    1906 => "10000100",
    1907 => "10000100",
    1908 => "10000100",
    1909 => "10000100",
    1910 => "10000100",
    1911 => "10000100",
    1912 => "10000100",
    1913 => "10000100",
    1914 => "10000100",
    1915 => "10000100",
    1916 => "10000100",
    1917 => "10000100",
    1918 => "10000100",
    1919 => "10000100",
    1920 => "10000100",
    1921 => "10000100",
    1922 => "10000011",
    1923 => "10000011",
    1924 => "10000011",
    1925 => "10000011",
    1926 => "10000011",
    1927 => "10000011",
    1928 => "10000011",
    1929 => "10000011",
    1930 => "10000011",
    1931 => "10000011",
    1932 => "10000011",
    1933 => "10000011",
    1934 => "10000011",
    1935 => "10000011",
    1936 => "10000011",
    1937 => "10000011",
    1938 => "10000011",
    1939 => "10000011",
    1940 => "10000011",
    1941 => "10000011",
    1942 => "10000011",
    1943 => "10000011",
    1944 => "10000011",
    1945 => "10000011",
    1946 => "10000011",
    1947 => "10000011",
    1948 => "10000011",
    1949 => "10000011",
    1950 => "10000011",
    1951 => "10000011",
    1952 => "10000011",
    1953 => "10000011",
    1954 => "10000010",
    1955 => "10000010",
    1956 => "10000010",
    1957 => "10000010",
    1958 => "10000010",
    1959 => "10000010",
    1960 => "10000010",
    1961 => "10000010",
    1962 => "10000010",
    1963 => "10000010",
    1964 => "10000010",
    1965 => "10000010",
    1966 => "10000010",
    1967 => "10000010",
    1968 => "10000010",
    1969 => "10000010",
    1970 => "10000010",
    1971 => "10000010",
    1972 => "10000010",
    1973 => "10000010",
    1974 => "10000010",
    1975 => "10000010",
    1976 => "10000010",
    1977 => "10000010",
    1978 => "10000010",
    1979 => "10000010",
    1980 => "10000010",
    1981 => "10000010",
    1982 => "10000010",
    1983 => "10000010",
    1984 => "10000010",
    1985 => "10000001",
    1986 => "10000001",
    1987 => "10000001",
    1988 => "10000001",
    1989 => "10000001",
    1990 => "10000001",
    1991 => "10000001",
    1992 => "10000001",
    1993 => "10000001",
    1994 => "10000001",
    1995 => "10000001",
    1996 => "10000001",
    1997 => "10000001",
    1998 => "10000001",
    1999 => "10000001",
    2000 => "10000001",
    2001 => "10000001",
    2002 => "10000001",
    2003 => "10000001",
    2004 => "10000001",
    2005 => "10000001",
    2006 => "10000001",
    2007 => "10000001",
    2008 => "10000001",
    2009 => "10000001",
    2010 => "10000001",
    2011 => "10000001",
    2012 => "10000001",
    2013 => "10000001",
    2014 => "10000001",
    2015 => "10000001",
    2016 => "10000001",
    2017 => "10000000",
    2018 => "10000000",
    2019 => "10000000",
    2020 => "10000000",
    2021 => "10000000",
    2022 => "10000000",
    2023 => "10000000",
    2024 => "10000000",
    2025 => "10000000",
    2026 => "10000000",
    2027 => "10000000",
    2028 => "10000000",
    2029 => "10000000",
    2030 => "10000000",
    2031 => "10000000",
    2032 => "10000000",
    2033 => "10000000",
    2034 => "10000000",
    2035 => "10000000",
    2036 => "10000000",
    2037 => "10000000",
    2038 => "10000000",
    2039 => "10000000",
    2040 => "10000000",
    2041 => "10000000",
    2042 => "10000000",
    2043 => "10000000",
    2044 => "10000000",
    2045 => "10000000",
    2046 => "10000000",
    2047 => "10000000",
    2048 => "01111111",
    2049 => "01111111",
    2050 => "01111111",
    2051 => "01111111",
    2052 => "01111111",
    2053 => "01111111",
    2054 => "01111111",
    2055 => "01111111",
    2056 => "01111111",
    2057 => "01111111",
    2058 => "01111111",
    2059 => "01111111",
    2060 => "01111111",
    2061 => "01111111",
    2062 => "01111111",
    2063 => "01111111",
    2064 => "01111111",
    2065 => "01111111",
    2066 => "01111111",
    2067 => "01111111",
    2068 => "01111111",
    2069 => "01111111",
    2070 => "01111111",
    2071 => "01111111",
    2072 => "01111111",
    2073 => "01111111",
    2074 => "01111111",
    2075 => "01111111",
    2076 => "01111111",
    2077 => "01111111",
    2078 => "01111111",
    2079 => "01111111",
    2080 => "01111111",
    2081 => "01111110",
    2082 => "01111110",
    2083 => "01111110",
    2084 => "01111110",
    2085 => "01111110",
    2086 => "01111110",
    2087 => "01111110",
    2088 => "01111110",
    2089 => "01111110",
    2090 => "01111110",
    2091 => "01111110",
    2092 => "01111110",
    2093 => "01111110",
    2094 => "01111110",
    2095 => "01111110",
    2096 => "01111110",
    2097 => "01111110",
    2098 => "01111110",
    2099 => "01111110",
    2100 => "01111110",
    2101 => "01111110",
    2102 => "01111110",
    2103 => "01111110",
    2104 => "01111110",
    2105 => "01111110",
    2106 => "01111110",
    2107 => "01111110",
    2108 => "01111110",
    2109 => "01111110",
    2110 => "01111110",
    2111 => "01111110",
    2112 => "01111110",
    2113 => "01111101",
    2114 => "01111101",
    2115 => "01111101",
    2116 => "01111101",
    2117 => "01111101",
    2118 => "01111101",
    2119 => "01111101",
    2120 => "01111101",
    2121 => "01111101",
    2122 => "01111101",
    2123 => "01111101",
    2124 => "01111101",
    2125 => "01111101",
    2126 => "01111101",
    2127 => "01111101",
    2128 => "01111101",
    2129 => "01111101",
    2130 => "01111101",
    2131 => "01111101",
    2132 => "01111101",
    2133 => "01111101",
    2134 => "01111101",
    2135 => "01111101",
    2136 => "01111101",
    2137 => "01111101",
    2138 => "01111101",
    2139 => "01111101",
    2140 => "01111101",
    2141 => "01111101",
    2142 => "01111101",
    2143 => "01111101",
    2144 => "01111101",
    2145 => "01111101",
    2146 => "01111100",
    2147 => "01111100",
    2148 => "01111100",
    2149 => "01111100",
    2150 => "01111100",
    2151 => "01111100",
    2152 => "01111100",
    2153 => "01111100",
    2154 => "01111100",
    2155 => "01111100",
    2156 => "01111100",
    2157 => "01111100",
    2158 => "01111100",
    2159 => "01111100",
    2160 => "01111100",
    2161 => "01111100",
    2162 => "01111100",
    2163 => "01111100",
    2164 => "01111100",
    2165 => "01111100",
    2166 => "01111100",
    2167 => "01111100",
    2168 => "01111100",
    2169 => "01111100",
    2170 => "01111100",
    2171 => "01111100",
    2172 => "01111100",
    2173 => "01111100",
    2174 => "01111100",
    2175 => "01111100",
    2176 => "01111100",
    2177 => "01111100",
    2178 => "01111011",
    2179 => "01111011",
    2180 => "01111011",
    2181 => "01111011",
    2182 => "01111011",
    2183 => "01111011",
    2184 => "01111011",
    2185 => "01111011",
    2186 => "01111011",
    2187 => "01111011",
    2188 => "01111011",
    2189 => "01111011",
    2190 => "01111011",
    2191 => "01111011",
    2192 => "01111011",
    2193 => "01111011",
    2194 => "01111011",
    2195 => "01111011",
    2196 => "01111011",
    2197 => "01111011",
    2198 => "01111011",
    2199 => "01111011",
    2200 => "01111011",
    2201 => "01111011",
    2202 => "01111011",
    2203 => "01111011",
    2204 => "01111011",
    2205 => "01111011",
    2206 => "01111011",
    2207 => "01111011",
    2208 => "01111011",
    2209 => "01111011",
    2210 => "01111011",
    2211 => "01111011",
    2212 => "01111010",
    2213 => "01111010",
    2214 => "01111010",
    2215 => "01111010",
    2216 => "01111010",
    2217 => "01111010",
    2218 => "01111010",
    2219 => "01111010",
    2220 => "01111010",
    2221 => "01111010",
    2222 => "01111010",
    2223 => "01111010",
    2224 => "01111010",
    2225 => "01111010",
    2226 => "01111010",
    2227 => "01111010",
    2228 => "01111010",
    2229 => "01111010",
    2230 => "01111010",
    2231 => "01111010",
    2232 => "01111010",
    2233 => "01111010",
    2234 => "01111010",
    2235 => "01111010",
    2236 => "01111010",
    2237 => "01111010",
    2238 => "01111010",
    2239 => "01111010",
    2240 => "01111010",
    2241 => "01111010",
    2242 => "01111010",
    2243 => "01111010",
    2244 => "01111010",
    2245 => "01111001",
    2246 => "01111001",
    2247 => "01111001",
    2248 => "01111001",
    2249 => "01111001",
    2250 => "01111001",
    2251 => "01111001",
    2252 => "01111001",
    2253 => "01111001",
    2254 => "01111001",
    2255 => "01111001",
    2256 => "01111001",
    2257 => "01111001",
    2258 => "01111001",
    2259 => "01111001",
    2260 => "01111001",
    2261 => "01111001",
    2262 => "01111001",
    2263 => "01111001",
    2264 => "01111001",
    2265 => "01111001",
    2266 => "01111001",
    2267 => "01111001",
    2268 => "01111001",
    2269 => "01111001",
    2270 => "01111001",
    2271 => "01111001",
    2272 => "01111001",
    2273 => "01111001",
    2274 => "01111001",
    2275 => "01111001",
    2276 => "01111001",
    2277 => "01111001",
    2278 => "01111001",
    2279 => "01111000",
    2280 => "01111000",
    2281 => "01111000",
    2282 => "01111000",
    2283 => "01111000",
    2284 => "01111000",
    2285 => "01111000",
    2286 => "01111000",
    2287 => "01111000",
    2288 => "01111000",
    2289 => "01111000",
    2290 => "01111000",
    2291 => "01111000",
    2292 => "01111000",
    2293 => "01111000",
    2294 => "01111000",
    2295 => "01111000",
    2296 => "01111000",
    2297 => "01111000",
    2298 => "01111000",
    2299 => "01111000",
    2300 => "01111000",
    2301 => "01111000",
    2302 => "01111000",
    2303 => "01111000",
    2304 => "01111000",
    2305 => "01111000",
    2306 => "01111000",
    2307 => "01111000",
    2308 => "01111000",
    2309 => "01111000",
    2310 => "01111000",
    2311 => "01111000",
    2312 => "01110111",
    2313 => "01110111",
    2314 => "01110111",
    2315 => "01110111",
    2316 => "01110111",
    2317 => "01110111",
    2318 => "01110111",
    2319 => "01110111",
    2320 => "01110111",
    2321 => "01110111",
    2322 => "01110111",
    2323 => "01110111",
    2324 => "01110111",
    2325 => "01110111",
    2326 => "01110111",
    2327 => "01110111",
    2328 => "01110111",
    2329 => "01110111",
    2330 => "01110111",
    2331 => "01110111",
    2332 => "01110111",
    2333 => "01110111",
    2334 => "01110111",
    2335 => "01110111",
    2336 => "01110111",
    2337 => "01110111",
    2338 => "01110111",
    2339 => "01110111",
    2340 => "01110111",
    2341 => "01110111",
    2342 => "01110111",
    2343 => "01110111",
    2344 => "01110111",
    2345 => "01110111",
    2346 => "01110111",
    2347 => "01110110",
    2348 => "01110110",
    2349 => "01110110",
    2350 => "01110110",
    2351 => "01110110",
    2352 => "01110110",
    2353 => "01110110",
    2354 => "01110110",
    2355 => "01110110",
    2356 => "01110110",
    2357 => "01110110",
    2358 => "01110110",
    2359 => "01110110",
    2360 => "01110110",
    2361 => "01110110",
    2362 => "01110110",
    2363 => "01110110",
    2364 => "01110110",
    2365 => "01110110",
    2366 => "01110110",
    2367 => "01110110",
    2368 => "01110110",
    2369 => "01110110",
    2370 => "01110110",
    2371 => "01110110",
    2372 => "01110110",
    2373 => "01110110",
    2374 => "01110110",
    2375 => "01110110",
    2376 => "01110110",
    2377 => "01110110",
    2378 => "01110110",
    2379 => "01110110",
    2380 => "01110110",
    2381 => "01110101",
    2382 => "01110101",
    2383 => "01110101",
    2384 => "01110101",
    2385 => "01110101",
    2386 => "01110101",
    2387 => "01110101",
    2388 => "01110101",
    2389 => "01110101",
    2390 => "01110101",
    2391 => "01110101",
    2392 => "01110101",
    2393 => "01110101",
    2394 => "01110101",
    2395 => "01110101",
    2396 => "01110101",
    2397 => "01110101",
    2398 => "01110101",
    2399 => "01110101",
    2400 => "01110101",
    2401 => "01110101",
    2402 => "01110101",
    2403 => "01110101",
    2404 => "01110101",
    2405 => "01110101",
    2406 => "01110101",
    2407 => "01110101",
    2408 => "01110101",
    2409 => "01110101",
    2410 => "01110101",
    2411 => "01110101",
    2412 => "01110101",
    2413 => "01110101",
    2414 => "01110101",
    2415 => "01110101",
    2416 => "01110100",
    2417 => "01110100",
    2418 => "01110100",
    2419 => "01110100",
    2420 => "01110100",
    2421 => "01110100",
    2422 => "01110100",
    2423 => "01110100",
    2424 => "01110100",
    2425 => "01110100",
    2426 => "01110100",
    2427 => "01110100",
    2428 => "01110100",
    2429 => "01110100",
    2430 => "01110100",
    2431 => "01110100",
    2432 => "01110100",
    2433 => "01110100",
    2434 => "01110100",
    2435 => "01110100",
    2436 => "01110100",
    2437 => "01110100",
    2438 => "01110100",
    2439 => "01110100",
    2440 => "01110100",
    2441 => "01110100",
    2442 => "01110100",
    2443 => "01110100",
    2444 => "01110100",
    2445 => "01110100",
    2446 => "01110100",
    2447 => "01110100",
    2448 => "01110100",
    2449 => "01110100",
    2450 => "01110011",
    2451 => "01110011",
    2452 => "01110011",
    2453 => "01110011",
    2454 => "01110011",
    2455 => "01110011",
    2456 => "01110011",
    2457 => "01110011",
    2458 => "01110011",
    2459 => "01110011",
    2460 => "01110011",
    2461 => "01110011",
    2462 => "01110011",
    2463 => "01110011",
    2464 => "01110011",
    2465 => "01110011",
    2466 => "01110011",
    2467 => "01110011",
    2468 => "01110011",
    2469 => "01110011",
    2470 => "01110011",
    2471 => "01110011",
    2472 => "01110011",
    2473 => "01110011",
    2474 => "01110011",
    2475 => "01110011",
    2476 => "01110011",
    2477 => "01110011",
    2478 => "01110011",
    2479 => "01110011",
    2480 => "01110011",
    2481 => "01110011",
    2482 => "01110011",
    2483 => "01110011",
    2484 => "01110011",
    2485 => "01110011",
    2486 => "01110010",
    2487 => "01110010",
    2488 => "01110010",
    2489 => "01110010",
    2490 => "01110010",
    2491 => "01110010",
    2492 => "01110010",
    2493 => "01110010",
    2494 => "01110010",
    2495 => "01110010",
    2496 => "01110010",
    2497 => "01110010",
    2498 => "01110010",
    2499 => "01110010",
    2500 => "01110010",
    2501 => "01110010",
    2502 => "01110010",
    2503 => "01110010",
    2504 => "01110010",
    2505 => "01110010",
    2506 => "01110010",
    2507 => "01110010",
    2508 => "01110010",
    2509 => "01110010",
    2510 => "01110010",
    2511 => "01110010",
    2512 => "01110010",
    2513 => "01110010",
    2514 => "01110010",
    2515 => "01110010",
    2516 => "01110010",
    2517 => "01110010",
    2518 => "01110010",
    2519 => "01110010",
    2520 => "01110010",
    2521 => "01110001",
    2522 => "01110001",
    2523 => "01110001",
    2524 => "01110001",
    2525 => "01110001",
    2526 => "01110001",
    2527 => "01110001",
    2528 => "01110001",
    2529 => "01110001",
    2530 => "01110001",
    2531 => "01110001",
    2532 => "01110001",
    2533 => "01110001",
    2534 => "01110001",
    2535 => "01110001",
    2536 => "01110001",
    2537 => "01110001",
    2538 => "01110001",
    2539 => "01110001",
    2540 => "01110001",
    2541 => "01110001",
    2542 => "01110001",
    2543 => "01110001",
    2544 => "01110001",
    2545 => "01110001",
    2546 => "01110001",
    2547 => "01110001",
    2548 => "01110001",
    2549 => "01110001",
    2550 => "01110001",
    2551 => "01110001",
    2552 => "01110001",
    2553 => "01110001",
    2554 => "01110001",
    2555 => "01110001",
    2556 => "01110001",
    2557 => "01110000",
    2558 => "01110000",
    2559 => "01110000",
    2560 => "01110000",
    2561 => "01110000",
    2562 => "01110000",
    2563 => "01110000",
    2564 => "01110000",
    2565 => "01110000",
    2566 => "01110000",
    2567 => "01110000",
    2568 => "01110000",
    2569 => "01110000",
    2570 => "01110000",
    2571 => "01110000",
    2572 => "01110000",
    2573 => "01110000",
    2574 => "01110000",
    2575 => "01110000",
    2576 => "01110000",
    2577 => "01110000",
    2578 => "01110000",
    2579 => "01110000",
    2580 => "01110000",
    2581 => "01110000",
    2582 => "01110000",
    2583 => "01110000",
    2584 => "01110000",
    2585 => "01110000",
    2586 => "01110000",
    2587 => "01110000",
    2588 => "01110000",
    2589 => "01110000",
    2590 => "01110000",
    2591 => "01110000",
    2592 => "01101111",
    2593 => "01101111",
    2594 => "01101111",
    2595 => "01101111",
    2596 => "01101111",
    2597 => "01101111",
    2598 => "01101111",
    2599 => "01101111",
    2600 => "01101111",
    2601 => "01101111",
    2602 => "01101111",
    2603 => "01101111",
    2604 => "01101111",
    2605 => "01101111",
    2606 => "01101111",
    2607 => "01101111",
    2608 => "01101111",
    2609 => "01101111",
    2610 => "01101111",
    2611 => "01101111",
    2612 => "01101111",
    2613 => "01101111",
    2614 => "01101111",
    2615 => "01101111",
    2616 => "01101111",
    2617 => "01101111",
    2618 => "01101111",
    2619 => "01101111",
    2620 => "01101111",
    2621 => "01101111",
    2622 => "01101111",
    2623 => "01101111",
    2624 => "01101111",
    2625 => "01101111",
    2626 => "01101111",
    2627 => "01101111",
    2628 => "01101111",
    2629 => "01101110",
    2630 => "01101110",
    2631 => "01101110",
    2632 => "01101110",
    2633 => "01101110",
    2634 => "01101110",
    2635 => "01101110",
    2636 => "01101110",
    2637 => "01101110",
    2638 => "01101110",
    2639 => "01101110",
    2640 => "01101110",
    2641 => "01101110",
    2642 => "01101110",
    2643 => "01101110",
    2644 => "01101110",
    2645 => "01101110",
    2646 => "01101110",
    2647 => "01101110",
    2648 => "01101110",
    2649 => "01101110",
    2650 => "01101110",
    2651 => "01101110",
    2652 => "01101110",
    2653 => "01101110",
    2654 => "01101110",
    2655 => "01101110",
    2656 => "01101110",
    2657 => "01101110",
    2658 => "01101110",
    2659 => "01101110",
    2660 => "01101110",
    2661 => "01101110",
    2662 => "01101110",
    2663 => "01101110",
    2664 => "01101110",
    2665 => "01101101",
    2666 => "01101101",
    2667 => "01101101",
    2668 => "01101101",
    2669 => "01101101",
    2670 => "01101101",
    2671 => "01101101",
    2672 => "01101101",
    2673 => "01101101",
    2674 => "01101101",
    2675 => "01101101",
    2676 => "01101101",
    2677 => "01101101",
    2678 => "01101101",
    2679 => "01101101",
    2680 => "01101101",
    2681 => "01101101",
    2682 => "01101101",
    2683 => "01101101",
    2684 => "01101101",
    2685 => "01101101",
    2686 => "01101101",
    2687 => "01101101",
    2688 => "01101101",
    2689 => "01101101",
    2690 => "01101101",
    2691 => "01101101",
    2692 => "01101101",
    2693 => "01101101",
    2694 => "01101101",
    2695 => "01101101",
    2696 => "01101101",
    2697 => "01101101",
    2698 => "01101101",
    2699 => "01101101",
    2700 => "01101101",
    2701 => "01101101",
    2702 => "01101100",
    2703 => "01101100",
    2704 => "01101100",
    2705 => "01101100",
    2706 => "01101100",
    2707 => "01101100",
    2708 => "01101100",
    2709 => "01101100",
    2710 => "01101100",
    2711 => "01101100",
    2712 => "01101100",
    2713 => "01101100",
    2714 => "01101100",
    2715 => "01101100",
    2716 => "01101100",
    2717 => "01101100",
    2718 => "01101100",
    2719 => "01101100",
    2720 => "01101100",
    2721 => "01101100",
    2722 => "01101100",
    2723 => "01101100",
    2724 => "01101100",
    2725 => "01101100",
    2726 => "01101100",
    2727 => "01101100",
    2728 => "01101100",
    2729 => "01101100",
    2730 => "01101100",
    2731 => "01101100",
    2732 => "01101100",
    2733 => "01101100",
    2734 => "01101100",
    2735 => "01101100",
    2736 => "01101100",
    2737 => "01101100",
    2738 => "01101011",
    2739 => "01101011",
    2740 => "01101011",
    2741 => "01101011",
    2742 => "01101011",
    2743 => "01101011",
    2744 => "01101011",
    2745 => "01101011",
    2746 => "01101011",
    2747 => "01101011",
    2748 => "01101011",
    2749 => "01101011",
    2750 => "01101011",
    2751 => "01101011",
    2752 => "01101011",
    2753 => "01101011",
    2754 => "01101011",
    2755 => "01101011",
    2756 => "01101011",
    2757 => "01101011",
    2758 => "01101011",
    2759 => "01101011",
    2760 => "01101011",
    2761 => "01101011",
    2762 => "01101011",
    2763 => "01101011",
    2764 => "01101011",
    2765 => "01101011",
    2766 => "01101011",
    2767 => "01101011",
    2768 => "01101011",
    2769 => "01101011",
    2770 => "01101011",
    2771 => "01101011",
    2772 => "01101011",
    2773 => "01101011",
    2774 => "01101011",
    2775 => "01101011",
    2776 => "01101010",
    2777 => "01101010",
    2778 => "01101010",
    2779 => "01101010",
    2780 => "01101010",
    2781 => "01101010",
    2782 => "01101010",
    2783 => "01101010",
    2784 => "01101010",
    2785 => "01101010",
    2786 => "01101010",
    2787 => "01101010",
    2788 => "01101010",
    2789 => "01101010",
    2790 => "01101010",
    2791 => "01101010",
    2792 => "01101010",
    2793 => "01101010",
    2794 => "01101010",
    2795 => "01101010",
    2796 => "01101010",
    2797 => "01101010",
    2798 => "01101010",
    2799 => "01101010",
    2800 => "01101010",
    2801 => "01101010",
    2802 => "01101010",
    2803 => "01101010",
    2804 => "01101010",
    2805 => "01101010",
    2806 => "01101010",
    2807 => "01101010",
    2808 => "01101010",
    2809 => "01101010",
    2810 => "01101010",
    2811 => "01101010",
    2812 => "01101010",
    2813 => "01101001",
    2814 => "01101001",
    2815 => "01101001",
    2816 => "01101001",
    2817 => "01101001",
    2818 => "01101001",
    2819 => "01101001",
    2820 => "01101001",
    2821 => "01101001",
    2822 => "01101001",
    2823 => "01101001",
    2824 => "01101001",
    2825 => "01101001",
    2826 => "01101001",
    2827 => "01101001",
    2828 => "01101001",
    2829 => "01101001",
    2830 => "01101001",
    2831 => "01101001",
    2832 => "01101001",
    2833 => "01101001",
    2834 => "01101001",
    2835 => "01101001",
    2836 => "01101001",
    2837 => "01101001",
    2838 => "01101001",
    2839 => "01101001",
    2840 => "01101001",
    2841 => "01101001",
    2842 => "01101001",
    2843 => "01101001",
    2844 => "01101001",
    2845 => "01101001",
    2846 => "01101001",
    2847 => "01101001",
    2848 => "01101001",
    2849 => "01101001",
    2850 => "01101001",
    2851 => "01101000",
    2852 => "01101000",
    2853 => "01101000",
    2854 => "01101000",
    2855 => "01101000",
    2856 => "01101000",
    2857 => "01101000",
    2858 => "01101000",
    2859 => "01101000",
    2860 => "01101000",
    2861 => "01101000",
    2862 => "01101000",
    2863 => "01101000",
    2864 => "01101000",
    2865 => "01101000",
    2866 => "01101000",
    2867 => "01101000",
    2868 => "01101000",
    2869 => "01101000",
    2870 => "01101000",
    2871 => "01101000",
    2872 => "01101000",
    2873 => "01101000",
    2874 => "01101000",
    2875 => "01101000",
    2876 => "01101000",
    2877 => "01101000",
    2878 => "01101000",
    2879 => "01101000",
    2880 => "01101000",
    2881 => "01101000",
    2882 => "01101000",
    2883 => "01101000",
    2884 => "01101000",
    2885 => "01101000",
    2886 => "01101000",
    2887 => "01101000",
    2888 => "01100111",
    2889 => "01100111",
    2890 => "01100111",
    2891 => "01100111",
    2892 => "01100111",
    2893 => "01100111",
    2894 => "01100111",
    2895 => "01100111",
    2896 => "01100111",
    2897 => "01100111",
    2898 => "01100111",
    2899 => "01100111",
    2900 => "01100111",
    2901 => "01100111",
    2902 => "01100111",
    2903 => "01100111",
    2904 => "01100111",
    2905 => "01100111",
    2906 => "01100111",
    2907 => "01100111",
    2908 => "01100111",
    2909 => "01100111",
    2910 => "01100111",
    2911 => "01100111",
    2912 => "01100111",
    2913 => "01100111",
    2914 => "01100111",
    2915 => "01100111",
    2916 => "01100111",
    2917 => "01100111",
    2918 => "01100111",
    2919 => "01100111",
    2920 => "01100111",
    2921 => "01100111",
    2922 => "01100111",
    2923 => "01100111",
    2924 => "01100111",
    2925 => "01100111",
    2926 => "01100111",
    2927 => "01100110",
    2928 => "01100110",
    2929 => "01100110",
    2930 => "01100110",
    2931 => "01100110",
    2932 => "01100110",
    2933 => "01100110",
    2934 => "01100110",
    2935 => "01100110",
    2936 => "01100110",
    2937 => "01100110",
    2938 => "01100110",
    2939 => "01100110",
    2940 => "01100110",
    2941 => "01100110",
    2942 => "01100110",
    2943 => "01100110",
    2944 => "01100110",
    2945 => "01100110",
    2946 => "01100110",
    2947 => "01100110",
    2948 => "01100110",
    2949 => "01100110",
    2950 => "01100110",
    2951 => "01100110",
    2952 => "01100110",
    2953 => "01100110",
    2954 => "01100110",
    2955 => "01100110",
    2956 => "01100110",
    2957 => "01100110",
    2958 => "01100110",
    2959 => "01100110",
    2960 => "01100110",
    2961 => "01100110",
    2962 => "01100110",
    2963 => "01100110",
    2964 => "01100110",
    2965 => "01100101",
    2966 => "01100101",
    2967 => "01100101",
    2968 => "01100101",
    2969 => "01100101",
    2970 => "01100101",
    2971 => "01100101",
    2972 => "01100101",
    2973 => "01100101",
    2974 => "01100101",
    2975 => "01100101",
    2976 => "01100101",
    2977 => "01100101",
    2978 => "01100101",
    2979 => "01100101",
    2980 => "01100101",
    2981 => "01100101",
    2982 => "01100101",
    2983 => "01100101",
    2984 => "01100101",
    2985 => "01100101",
    2986 => "01100101",
    2987 => "01100101",
    2988 => "01100101",
    2989 => "01100101",
    2990 => "01100101",
    2991 => "01100101",
    2992 => "01100101",
    2993 => "01100101",
    2994 => "01100101",
    2995 => "01100101",
    2996 => "01100101",
    2997 => "01100101",
    2998 => "01100101",
    2999 => "01100101",
    3000 => "01100101",
    3001 => "01100101",
    3002 => "01100101",
    3003 => "01100101",
    3004 => "01100100",
    3005 => "01100100",
    3006 => "01100100",
    3007 => "01100100",
    3008 => "01100100",
    3009 => "01100100",
    3010 => "01100100",
    3011 => "01100100",
    3012 => "01100100",
    3013 => "01100100",
    3014 => "01100100",
    3015 => "01100100",
    3016 => "01100100",
    3017 => "01100100",
    3018 => "01100100",
    3019 => "01100100",
    3020 => "01100100",
    3021 => "01100100",
    3022 => "01100100",
    3023 => "01100100",
    3024 => "01100100",
    3025 => "01100100",
    3026 => "01100100",
    3027 => "01100100",
    3028 => "01100100",
    3029 => "01100100",
    3030 => "01100100",
    3031 => "01100100",
    3032 => "01100100",
    3033 => "01100100",
    3034 => "01100100",
    3035 => "01100100",
    3036 => "01100100",
    3037 => "01100100",
    3038 => "01100100",
    3039 => "01100100",
    3040 => "01100100",
    3041 => "01100100",
    3042 => "01100011",
    3043 => "01100011",
    3044 => "01100011",
    3045 => "01100011",
    3046 => "01100011",
    3047 => "01100011",
    3048 => "01100011",
    3049 => "01100011",
    3050 => "01100011",
    3051 => "01100011",
    3052 => "01100011",
    3053 => "01100011",
    3054 => "01100011",
    3055 => "01100011",
    3056 => "01100011",
    3057 => "01100011",
    3058 => "01100011",
    3059 => "01100011",
    3060 => "01100011",
    3061 => "01100011",
    3062 => "01100011",
    3063 => "01100011",
    3064 => "01100011",
    3065 => "01100011",
    3066 => "01100011",
    3067 => "01100011",
    3068 => "01100011",
    3069 => "01100011",
    3070 => "01100011",
    3071 => "01100011",
    3072 => "01100011",
    3073 => "01100011",
    3074 => "01100011",
    3075 => "01100011",
    3076 => "01100011",
    3077 => "01100011",
    3078 => "01100011",
    3079 => "01100011",
    3080 => "01100011",
    3081 => "01100011",
    3082 => "01100010",
    3083 => "01100010",
    3084 => "01100010",
    3085 => "01100010",
    3086 => "01100010",
    3087 => "01100010",
    3088 => "01100010",
    3089 => "01100010",
    3090 => "01100010",
    3091 => "01100010",
    3092 => "01100010",
    3093 => "01100010",
    3094 => "01100010",
    3095 => "01100010",
    3096 => "01100010",
    3097 => "01100010",
    3098 => "01100010",
    3099 => "01100010",
    3100 => "01100010",
    3101 => "01100010",
    3102 => "01100010",
    3103 => "01100010",
    3104 => "01100010",
    3105 => "01100010",
    3106 => "01100010",
    3107 => "01100010",
    3108 => "01100010",
    3109 => "01100010",
    3110 => "01100010",
    3111 => "01100010",
    3112 => "01100010",
    3113 => "01100010",
    3114 => "01100010",
    3115 => "01100010",
    3116 => "01100010",
    3117 => "01100010",
    3118 => "01100010",
    3119 => "01100010",
    3120 => "01100010",
    3121 => "01100001",
    3122 => "01100001",
    3123 => "01100001",
    3124 => "01100001",
    3125 => "01100001",
    3126 => "01100001",
    3127 => "01100001",
    3128 => "01100001",
    3129 => "01100001",
    3130 => "01100001",
    3131 => "01100001",
    3132 => "01100001",
    3133 => "01100001",
    3134 => "01100001",
    3135 => "01100001",
    3136 => "01100001",
    3137 => "01100001",
    3138 => "01100001",
    3139 => "01100001",
    3140 => "01100001",
    3141 => "01100001",
    3142 => "01100001",
    3143 => "01100001",
    3144 => "01100001",
    3145 => "01100001",
    3146 => "01100001",
    3147 => "01100001",
    3148 => "01100001",
    3149 => "01100001",
    3150 => "01100001",
    3151 => "01100001",
    3152 => "01100001",
    3153 => "01100001",
    3154 => "01100001",
    3155 => "01100001",
    3156 => "01100001",
    3157 => "01100001",
    3158 => "01100001",
    3159 => "01100001",
    3160 => "01100001",
    3161 => "01100000",
    3162 => "01100000",
    3163 => "01100000",
    3164 => "01100000",
    3165 => "01100000",
    3166 => "01100000",
    3167 => "01100000",
    3168 => "01100000",
    3169 => "01100000",
    3170 => "01100000",
    3171 => "01100000",
    3172 => "01100000",
    3173 => "01100000",
    3174 => "01100000",
    3175 => "01100000",
    3176 => "01100000",
    3177 => "01100000",
    3178 => "01100000",
    3179 => "01100000",
    3180 => "01100000",
    3181 => "01100000",
    3182 => "01100000",
    3183 => "01100000",
    3184 => "01100000",
    3185 => "01100000",
    3186 => "01100000",
    3187 => "01100000",
    3188 => "01100000",
    3189 => "01100000",
    3190 => "01100000",
    3191 => "01100000",
    3192 => "01100000",
    3193 => "01100000",
    3194 => "01100000",
    3195 => "01100000",
    3196 => "01100000",
    3197 => "01100000",
    3198 => "01100000",
    3199 => "01100000",
    3200 => "01011111",
    3201 => "01011111",
    3202 => "01011111",
    3203 => "01011111",
    3204 => "01011111",
    3205 => "01011111",
    3206 => "01011111",
    3207 => "01011111",
    3208 => "01011111",
    3209 => "01011111",
    3210 => "01011111",
    3211 => "01011111",
    3212 => "01011111",
    3213 => "01011111",
    3214 => "01011111",
    3215 => "01011111",
    3216 => "01011111",
    3217 => "01011111",
    3218 => "01011111",
    3219 => "01011111",
    3220 => "01011111",
    3221 => "01011111",
    3222 => "01011111",
    3223 => "01011111",
    3224 => "01011111",
    3225 => "01011111",
    3226 => "01011111",
    3227 => "01011111",
    3228 => "01011111",
    3229 => "01011111",
    3230 => "01011111",
    3231 => "01011111",
    3232 => "01011111",
    3233 => "01011111",
    3234 => "01011111",
    3235 => "01011111",
    3236 => "01011111",
    3237 => "01011111",
    3238 => "01011111",
    3239 => "01011111",
    3240 => "01011111",
    3241 => "01011110",
    3242 => "01011110",
    3243 => "01011110",
    3244 => "01011110",
    3245 => "01011110",
    3246 => "01011110",
    3247 => "01011110",
    3248 => "01011110",
    3249 => "01011110",
    3250 => "01011110",
    3251 => "01011110",
    3252 => "01011110",
    3253 => "01011110",
    3254 => "01011110",
    3255 => "01011110",
    3256 => "01011110",
    3257 => "01011110",
    3258 => "01011110",
    3259 => "01011110",
    3260 => "01011110",
    3261 => "01011110",
    3262 => "01011110",
    3263 => "01011110",
    3264 => "01011110",
    3265 => "01011110",
    3266 => "01011110",
    3267 => "01011110",
    3268 => "01011110",
    3269 => "01011110",
    3270 => "01011110",
    3271 => "01011110",
    3272 => "01011110",
    3273 => "01011110",
    3274 => "01011110",
    3275 => "01011110",
    3276 => "01011110",
    3277 => "01011110",
    3278 => "01011110",
    3279 => "01011110",
    3280 => "01011110",
    3281 => "01011101",
    3282 => "01011101",
    3283 => "01011101",
    3284 => "01011101",
    3285 => "01011101",
    3286 => "01011101",
    3287 => "01011101",
    3288 => "01011101",
    3289 => "01011101",
    3290 => "01011101",
    3291 => "01011101",
    3292 => "01011101",
    3293 => "01011101",
    3294 => "01011101",
    3295 => "01011101",
    3296 => "01011101",
    3297 => "01011101",
    3298 => "01011101",
    3299 => "01011101",
    3300 => "01011101",
    3301 => "01011101",
    3302 => "01011101",
    3303 => "01011101",
    3304 => "01011101",
    3305 => "01011101",
    3306 => "01011101",
    3307 => "01011101",
    3308 => "01011101",
    3309 => "01011101",
    3310 => "01011101",
    3311 => "01011101",
    3312 => "01011101",
    3313 => "01011101",
    3314 => "01011101",
    3315 => "01011101",
    3316 => "01011101",
    3317 => "01011101",
    3318 => "01011101",
    3319 => "01011101",
    3320 => "01011101",
    3321 => "01011101",
    3322 => "01011100",
    3323 => "01011100",
    3324 => "01011100",
    3325 => "01011100",
    3326 => "01011100",
    3327 => "01011100",
    3328 => "01011100",
    3329 => "01011100",
    3330 => "01011100",
    3331 => "01011100",
    3332 => "01011100",
    3333 => "01011100",
    3334 => "01011100",
    3335 => "01011100",
    3336 => "01011100",
    3337 => "01011100",
    3338 => "01011100",
    3339 => "01011100",
    3340 => "01011100",
    3341 => "01011100",
    3342 => "01011100",
    3343 => "01011100",
    3344 => "01011100",
    3345 => "01011100",
    3346 => "01011100",
    3347 => "01011100",
    3348 => "01011100",
    3349 => "01011100",
    3350 => "01011100",
    3351 => "01011100",
    3352 => "01011100",
    3353 => "01011100",
    3354 => "01011100",
    3355 => "01011100",
    3356 => "01011100",
    3357 => "01011100",
    3358 => "01011100",
    3359 => "01011100",
    3360 => "01011100",
    3361 => "01011100",
    3362 => "01011011",
    3363 => "01011011",
    3364 => "01011011",
    3365 => "01011011",
    3366 => "01011011",
    3367 => "01011011",
    3368 => "01011011",
    3369 => "01011011",
    3370 => "01011011",
    3371 => "01011011",
    3372 => "01011011",
    3373 => "01011011",
    3374 => "01011011",
    3375 => "01011011",
    3376 => "01011011",
    3377 => "01011011",
    3378 => "01011011",
    3379 => "01011011",
    3380 => "01011011",
    3381 => "01011011",
    3382 => "01011011",
    3383 => "01011011",
    3384 => "01011011",
    3385 => "01011011",
    3386 => "01011011",
    3387 => "01011011",
    3388 => "01011011",
    3389 => "01011011",
    3390 => "01011011",
    3391 => "01011011",
    3392 => "01011011",
    3393 => "01011011",
    3394 => "01011011",
    3395 => "01011011",
    3396 => "01011011",
    3397 => "01011011",
    3398 => "01011011",
    3399 => "01011011",
    3400 => "01011011",
    3401 => "01011011",
    3402 => "01011011",
    3403 => "01011011",
    3404 => "01011010",
    3405 => "01011010",
    3406 => "01011010",
    3407 => "01011010",
    3408 => "01011010",
    3409 => "01011010",
    3410 => "01011010",
    3411 => "01011010",
    3412 => "01011010",
    3413 => "01011010",
    3414 => "01011010",
    3415 => "01011010",
    3416 => "01011010",
    3417 => "01011010",
    3418 => "01011010",
    3419 => "01011010",
    3420 => "01011010",
    3421 => "01011010",
    3422 => "01011010",
    3423 => "01011010",
    3424 => "01011010",
    3425 => "01011010",
    3426 => "01011010",
    3427 => "01011010",
    3428 => "01011010",
    3429 => "01011010",
    3430 => "01011010",
    3431 => "01011010",
    3432 => "01011010",
    3433 => "01011010",
    3434 => "01011010",
    3435 => "01011010",
    3436 => "01011010",
    3437 => "01011010",
    3438 => "01011010",
    3439 => "01011010",
    3440 => "01011010",
    3441 => "01011010",
    3442 => "01011010",
    3443 => "01011010",
    3444 => "01011010",
    3445 => "01011001",
    3446 => "01011001",
    3447 => "01011001",
    3448 => "01011001",
    3449 => "01011001",
    3450 => "01011001",
    3451 => "01011001",
    3452 => "01011001",
    3453 => "01011001",
    3454 => "01011001",
    3455 => "01011001",
    3456 => "01011001",
    3457 => "01011001",
    3458 => "01011001",
    3459 => "01011001",
    3460 => "01011001",
    3461 => "01011001",
    3462 => "01011001",
    3463 => "01011001",
    3464 => "01011001",
    3465 => "01011001",
    3466 => "01011001",
    3467 => "01011001",
    3468 => "01011001",
    3469 => "01011001",
    3470 => "01011001",
    3471 => "01011001",
    3472 => "01011001",
    3473 => "01011001",
    3474 => "01011001",
    3475 => "01011001",
    3476 => "01011001",
    3477 => "01011001",
    3478 => "01011001",
    3479 => "01011001",
    3480 => "01011001",
    3481 => "01011001",
    3482 => "01011001",
    3483 => "01011001",
    3484 => "01011001",
    3485 => "01011001",
    3486 => "01011001",
    3487 => "01011000",
    3488 => "01011000",
    3489 => "01011000",
    3490 => "01011000",
    3491 => "01011000",
    3492 => "01011000",
    3493 => "01011000",
    3494 => "01011000",
    3495 => "01011000",
    3496 => "01011000",
    3497 => "01011000",
    3498 => "01011000",
    3499 => "01011000",
    3500 => "01011000",
    3501 => "01011000",
    3502 => "01011000",
    3503 => "01011000",
    3504 => "01011000",
    3505 => "01011000",
    3506 => "01011000",
    3507 => "01011000",
    3508 => "01011000",
    3509 => "01011000",
    3510 => "01011000",
    3511 => "01011000",
    3512 => "01011000",
    3513 => "01011000",
    3514 => "01011000",
    3515 => "01011000",
    3516 => "01011000",
    3517 => "01011000",
    3518 => "01011000",
    3519 => "01011000",
    3520 => "01011000",
    3521 => "01011000",
    3522 => "01011000",
    3523 => "01011000",
    3524 => "01011000",
    3525 => "01011000",
    3526 => "01011000",
    3527 => "01011000",
    3528 => "01010111",
    3529 => "01010111",
    3530 => "01010111",
    3531 => "01010111",
    3532 => "01010111",
    3533 => "01010111",
    3534 => "01010111",
    3535 => "01010111",
    3536 => "01010111",
    3537 => "01010111",
    3538 => "01010111",
    3539 => "01010111",
    3540 => "01010111",
    3541 => "01010111",
    3542 => "01010111",
    3543 => "01010111",
    3544 => "01010111",
    3545 => "01010111",
    3546 => "01010111",
    3547 => "01010111",
    3548 => "01010111",
    3549 => "01010111",
    3550 => "01010111",
    3551 => "01010111",
    3552 => "01010111",
    3553 => "01010111",
    3554 => "01010111",
    3555 => "01010111",
    3556 => "01010111",
    3557 => "01010111",
    3558 => "01010111",
    3559 => "01010111",
    3560 => "01010111",
    3561 => "01010111",
    3562 => "01010111",
    3563 => "01010111",
    3564 => "01010111",
    3565 => "01010111",
    3566 => "01010111",
    3567 => "01010111",
    3568 => "01010111",
    3569 => "01010111",
    3570 => "01010111",
    3571 => "01010110",
    3572 => "01010110",
    3573 => "01010110",
    3574 => "01010110",
    3575 => "01010110",
    3576 => "01010110",
    3577 => "01010110",
    3578 => "01010110",
    3579 => "01010110",
    3580 => "01010110",
    3581 => "01010110",
    3582 => "01010110",
    3583 => "01010110",
    3584 => "01010110",
    3585 => "01010110",
    3586 => "01010110",
    3587 => "01010110",
    3588 => "01010110",
    3589 => "01010110",
    3590 => "01010110",
    3591 => "01010110",
    3592 => "01010110",
    3593 => "01010110",
    3594 => "01010110",
    3595 => "01010110",
    3596 => "01010110",
    3597 => "01010110",
    3598 => "01010110",
    3599 => "01010110",
    3600 => "01010110",
    3601 => "01010110",
    3602 => "01010110",
    3603 => "01010110",
    3604 => "01010110",
    3605 => "01010110",
    3606 => "01010110",
    3607 => "01010110",
    3608 => "01010110",
    3609 => "01010110",
    3610 => "01010110",
    3611 => "01010110",
    3612 => "01010110",
    3613 => "01010101",
    3614 => "01010101",
    3615 => "01010101",
    3616 => "01010101",
    3617 => "01010101",
    3618 => "01010101",
    3619 => "01010101",
    3620 => "01010101",
    3621 => "01010101",
    3622 => "01010101",
    3623 => "01010101",
    3624 => "01010101",
    3625 => "01010101",
    3626 => "01010101",
    3627 => "01010101",
    3628 => "01010101",
    3629 => "01010101",
    3630 => "01010101",
    3631 => "01010101",
    3632 => "01010101",
    3633 => "01010101",
    3634 => "01010101",
    3635 => "01010101",
    3636 => "01010101",
    3637 => "01010101",
    3638 => "01010101",
    3639 => "01010101",
    3640 => "01010101",
    3641 => "01010101",
    3642 => "01010101",
    3643 => "01010101",
    3644 => "01010101",
    3645 => "01010101",
    3646 => "01010101",
    3647 => "01010101",
    3648 => "01010101",
    3649 => "01010101",
    3650 => "01010101",
    3651 => "01010101",
    3652 => "01010101",
    3653 => "01010101",
    3654 => "01010101",
    3655 => "01010101",
    3656 => "01010100",
    3657 => "01010100",
    3658 => "01010100",
    3659 => "01010100",
    3660 => "01010100",
    3661 => "01010100",
    3662 => "01010100",
    3663 => "01010100",
    3664 => "01010100",
    3665 => "01010100",
    3666 => "01010100",
    3667 => "01010100",
    3668 => "01010100",
    3669 => "01010100",
    3670 => "01010100",
    3671 => "01010100",
    3672 => "01010100",
    3673 => "01010100",
    3674 => "01010100",
    3675 => "01010100",
    3676 => "01010100",
    3677 => "01010100",
    3678 => "01010100",
    3679 => "01010100",
    3680 => "01010100",
    3681 => "01010100",
    3682 => "01010100",
    3683 => "01010100",
    3684 => "01010100",
    3685 => "01010100",
    3686 => "01010100",
    3687 => "01010100",
    3688 => "01010100",
    3689 => "01010100",
    3690 => "01010100",
    3691 => "01010100",
    3692 => "01010100",
    3693 => "01010100",
    3694 => "01010100",
    3695 => "01010100",
    3696 => "01010100",
    3697 => "01010100",
    3698 => "01010011",
    3699 => "01010011",
    3700 => "01010011",
    3701 => "01010011",
    3702 => "01010011",
    3703 => "01010011",
    3704 => "01010011",
    3705 => "01010011",
    3706 => "01010011",
    3707 => "01010011",
    3708 => "01010011",
    3709 => "01010011",
    3710 => "01010011",
    3711 => "01010011",
    3712 => "01010011",
    3713 => "01010011",
    3714 => "01010011",
    3715 => "01010011",
    3716 => "01010011",
    3717 => "01010011",
    3718 => "01010011",
    3719 => "01010011",
    3720 => "01010011",
    3721 => "01010011",
    3722 => "01010011",
    3723 => "01010011",
    3724 => "01010011",
    3725 => "01010011",
    3726 => "01010011",
    3727 => "01010011",
    3728 => "01010011",
    3729 => "01010011",
    3730 => "01010011",
    3731 => "01010011",
    3732 => "01010011",
    3733 => "01010011",
    3734 => "01010011",
    3735 => "01010011",
    3736 => "01010011",
    3737 => "01010011",
    3738 => "01010011",
    3739 => "01010011",
    3740 => "01010011",
    3741 => "01010011",
    3742 => "01010010",
    3743 => "01010010",
    3744 => "01010010",
    3745 => "01010010",
    3746 => "01010010",
    3747 => "01010010",
    3748 => "01010010",
    3749 => "01010010",
    3750 => "01010010",
    3751 => "01010010",
    3752 => "01010010",
    3753 => "01010010",
    3754 => "01010010",
    3755 => "01010010",
    3756 => "01010010",
    3757 => "01010010",
    3758 => "01010010",
    3759 => "01010010",
    3760 => "01010010",
    3761 => "01010010",
    3762 => "01010010",
    3763 => "01010010",
    3764 => "01010010",
    3765 => "01010010",
    3766 => "01010010",
    3767 => "01010010",
    3768 => "01010010",
    3769 => "01010010",
    3770 => "01010010",
    3771 => "01010010",
    3772 => "01010010",
    3773 => "01010010",
    3774 => "01010010",
    3775 => "01010010",
    3776 => "01010010",
    3777 => "01010010",
    3778 => "01010010",
    3779 => "01010010",
    3780 => "01010010",
    3781 => "01010010",
    3782 => "01010010",
    3783 => "01010010",
    3784 => "01010010",
    3785 => "01010001",
    3786 => "01010001",
    3787 => "01010001",
    3788 => "01010001",
    3789 => "01010001",
    3790 => "01010001",
    3791 => "01010001",
    3792 => "01010001",
    3793 => "01010001",
    3794 => "01010001",
    3795 => "01010001",
    3796 => "01010001",
    3797 => "01010001",
    3798 => "01010001",
    3799 => "01010001",
    3800 => "01010001",
    3801 => "01010001",
    3802 => "01010001",
    3803 => "01010001",
    3804 => "01010001",
    3805 => "01010001",
    3806 => "01010001",
    3807 => "01010001",
    3808 => "01010001",
    3809 => "01010001",
    3810 => "01010001",
    3811 => "01010001",
    3812 => "01010001",
    3813 => "01010001",
    3814 => "01010001",
    3815 => "01010001",
    3816 => "01010001",
    3817 => "01010001",
    3818 => "01010001",
    3819 => "01010001",
    3820 => "01010001",
    3821 => "01010001",
    3822 => "01010001",
    3823 => "01010001",
    3824 => "01010001",
    3825 => "01010001",
    3826 => "01010001",
    3827 => "01010001",
    3828 => "01010001",
    3829 => "01010000",
    3830 => "01010000",
    3831 => "01010000",
    3832 => "01010000",
    3833 => "01010000",
    3834 => "01010000",
    3835 => "01010000",
    3836 => "01010000",
    3837 => "01010000",
    3838 => "01010000",
    3839 => "01010000",
    3840 => "01010000",
    3841 => "01010000",
    3842 => "01010000",
    3843 => "01010000",
    3844 => "01010000",
    3845 => "01010000",
    3846 => "01010000",
    3847 => "01010000",
    3848 => "01010000",
    3849 => "01010000",
    3850 => "01010000",
    3851 => "01010000",
    3852 => "01010000",
    3853 => "01010000",
    3854 => "01010000",
    3855 => "01010000",
    3856 => "01010000",
    3857 => "01010000",
    3858 => "01010000",
    3859 => "01010000",
    3860 => "01010000",
    3861 => "01010000",
    3862 => "01010000",
    3863 => "01010000",
    3864 => "01010000",
    3865 => "01010000",
    3866 => "01010000",
    3867 => "01010000",
    3868 => "01010000",
    3869 => "01010000",
    3870 => "01010000",
    3871 => "01010000",
    3872 => "01001111",
    3873 => "01001111",
    3874 => "01001111",
    3875 => "01001111",
    3876 => "01001111",
    3877 => "01001111",
    3878 => "01001111",
    3879 => "01001111",
    3880 => "01001111",
    3881 => "01001111",
    3882 => "01001111",
    3883 => "01001111",
    3884 => "01001111",
    3885 => "01001111",
    3886 => "01001111",
    3887 => "01001111",
    3888 => "01001111",
    3889 => "01001111",
    3890 => "01001111",
    3891 => "01001111",
    3892 => "01001111",
    3893 => "01001111",
    3894 => "01001111",
    3895 => "01001111",
    3896 => "01001111",
    3897 => "01001111",
    3898 => "01001111",
    3899 => "01001111",
    3900 => "01001111",
    3901 => "01001111",
    3902 => "01001111",
    3903 => "01001111",
    3904 => "01001111",
    3905 => "01001111",
    3906 => "01001111",
    3907 => "01001111",
    3908 => "01001111",
    3909 => "01001111",
    3910 => "01001111",
    3911 => "01001111",
    3912 => "01001111",
    3913 => "01001111",
    3914 => "01001111",
    3915 => "01001111",
    3916 => "01001111",
    3917 => "01001110",
    3918 => "01001110",
    3919 => "01001110",
    3920 => "01001110",
    3921 => "01001110",
    3922 => "01001110",
    3923 => "01001110",
    3924 => "01001110",
    3925 => "01001110",
    3926 => "01001110",
    3927 => "01001110",
    3928 => "01001110",
    3929 => "01001110",
    3930 => "01001110",
    3931 => "01001110",
    3932 => "01001110",
    3933 => "01001110",
    3934 => "01001110",
    3935 => "01001110",
    3936 => "01001110",
    3937 => "01001110",
    3938 => "01001110",
    3939 => "01001110",
    3940 => "01001110",
    3941 => "01001110",
    3942 => "01001110",
    3943 => "01001110",
    3944 => "01001110",
    3945 => "01001110",
    3946 => "01001110",
    3947 => "01001110",
    3948 => "01001110",
    3949 => "01001110",
    3950 => "01001110",
    3951 => "01001110",
    3952 => "01001110",
    3953 => "01001110",
    3954 => "01001110",
    3955 => "01001110",
    3956 => "01001110",
    3957 => "01001110",
    3958 => "01001110",
    3959 => "01001110",
    3960 => "01001110",
    3961 => "01001101",
    3962 => "01001101",
    3963 => "01001101",
    3964 => "01001101",
    3965 => "01001101",
    3966 => "01001101",
    3967 => "01001101",
    3968 => "01001101",
    3969 => "01001101",
    3970 => "01001101",
    3971 => "01001101",
    3972 => "01001101",
    3973 => "01001101",
    3974 => "01001101",
    3975 => "01001101",
    3976 => "01001101",
    3977 => "01001101",
    3978 => "01001101",
    3979 => "01001101",
    3980 => "01001101",
    3981 => "01001101",
    3982 => "01001101",
    3983 => "01001101",
    3984 => "01001101",
    3985 => "01001101",
    3986 => "01001101",
    3987 => "01001101",
    3988 => "01001101",
    3989 => "01001101",
    3990 => "01001101",
    3991 => "01001101",
    3992 => "01001101",
    3993 => "01001101",
    3994 => "01001101",
    3995 => "01001101",
    3996 => "01001101",
    3997 => "01001101",
    3998 => "01001101",
    3999 => "01001101",
    4000 => "01001101",
    4001 => "01001101",
    4002 => "01001101",
    4003 => "01001101",
    4004 => "01001101",
    4005 => "01001101",
    4006 => "01001100",
    4007 => "01001100",
    4008 => "01001100",
    4009 => "01001100",
    4010 => "01001100",
    4011 => "01001100",
    4012 => "01001100",
    4013 => "01001100",
    4014 => "01001100",
    4015 => "01001100",
    4016 => "01001100",
    4017 => "01001100",
    4018 => "01001100",
    4019 => "01001100",
    4020 => "01001100",
    4021 => "01001100",
    4022 => "01001100",
    4023 => "01001100",
    4024 => "01001100",
    4025 => "01001100",
    4026 => "01001100",
    4027 => "01001100",
    4028 => "01001100",
    4029 => "01001100",
    4030 => "01001100",
    4031 => "01001100",
    4032 => "01001100",
    4033 => "01001100",
    4034 => "01001100",
    4035 => "01001100",
    4036 => "01001100",
    4037 => "01001100",
    4038 => "01001100",
    4039 => "01001100",
    4040 => "01001100",
    4041 => "01001100",
    4042 => "01001100",
    4043 => "01001100",
    4044 => "01001100",
    4045 => "01001100",
    4046 => "01001100",
    4047 => "01001100",
    4048 => "01001100",
    4049 => "01001100",
    4050 => "01001011",
    4051 => "01001011",
    4052 => "01001011",
    4053 => "01001011",
    4054 => "01001011",
    4055 => "01001011",
    4056 => "01001011",
    4057 => "01001011",
    4058 => "01001011",
    4059 => "01001011",
    4060 => "01001011",
    4061 => "01001011",
    4062 => "01001011",
    4063 => "01001011",
    4064 => "01001011",
    4065 => "01001011",
    4066 => "01001011",
    4067 => "01001011",
    4068 => "01001011",
    4069 => "01001011",
    4070 => "01001011",
    4071 => "01001011",
    4072 => "01001011",
    4073 => "01001011",
    4074 => "01001011",
    4075 => "01001011",
    4076 => "01001011",
    4077 => "01001011",
    4078 => "01001011",
    4079 => "01001011",
    4080 => "01001011",
    4081 => "01001011",
    4082 => "01001011",
    4083 => "01001011",
    4084 => "01001011",
    4085 => "01001011",
    4086 => "01001011",
    4087 => "01001011",
    4088 => "01001011",
    4089 => "01001011",
    4090 => "01001011",
    4091 => "01001011",
    4092 => "01001011",
    4093 => "01001011",
    4094 => "01001011",
    4095 => "01001011",
    4096 => "01001010",
    4097 => "01001010",
    4098 => "01001010",
    4099 => "01001010",
    4100 => "01001010",
    4101 => "01001010",
    4102 => "01001010",
    4103 => "01001010",
    4104 => "01001010",
    4105 => "01001010",
    4106 => "01001010",
    4107 => "01001010",
    4108 => "01001010",
    4109 => "01001010",
    4110 => "01001010",
    4111 => "01001010",
    4112 => "01001010",
    4113 => "01001010",
    4114 => "01001010",
    4115 => "01001010",
    4116 => "01001010",
    4117 => "01001010",
    4118 => "01001010",
    4119 => "01001010",
    4120 => "01001010",
    4121 => "01001010",
    4122 => "01001010",
    4123 => "01001010",
    4124 => "01001010",
    4125 => "01001010",
    4126 => "01001010",
    4127 => "01001010",
    4128 => "01001010",
    4129 => "01001010",
    4130 => "01001010",
    4131 => "01001010",
    4132 => "01001010",
    4133 => "01001010",
    4134 => "01001010",
    4135 => "01001010",
    4136 => "01001010",
    4137 => "01001010",
    4138 => "01001010",
    4139 => "01001010",
    4140 => "01001010",
    4141 => "01001001",
    4142 => "01001001",
    4143 => "01001001",
    4144 => "01001001",
    4145 => "01001001",
    4146 => "01001001",
    4147 => "01001001",
    4148 => "01001001",
    4149 => "01001001",
    4150 => "01001001",
    4151 => "01001001",
    4152 => "01001001",
    4153 => "01001001",
    4154 => "01001001",
    4155 => "01001001",
    4156 => "01001001",
    4157 => "01001001",
    4158 => "01001001",
    4159 => "01001001",
    4160 => "01001001",
    4161 => "01001001",
    4162 => "01001001",
    4163 => "01001001",
    4164 => "01001001",
    4165 => "01001001",
    4166 => "01001001",
    4167 => "01001001",
    4168 => "01001001",
    4169 => "01001001",
    4170 => "01001001",
    4171 => "01001001",
    4172 => "01001001",
    4173 => "01001001",
    4174 => "01001001",
    4175 => "01001001",
    4176 => "01001001",
    4177 => "01001001",
    4178 => "01001001",
    4179 => "01001001",
    4180 => "01001001",
    4181 => "01001001",
    4182 => "01001001",
    4183 => "01001001",
    4184 => "01001001",
    4185 => "01001001",
    4186 => "01001001",
    4187 => "01001000",
    4188 => "01001000",
    4189 => "01001000",
    4190 => "01001000",
    4191 => "01001000",
    4192 => "01001000",
    4193 => "01001000",
    4194 => "01001000",
    4195 => "01001000",
    4196 => "01001000",
    4197 => "01001000",
    4198 => "01001000",
    4199 => "01001000",
    4200 => "01001000",
    4201 => "01001000",
    4202 => "01001000",
    4203 => "01001000",
    4204 => "01001000",
    4205 => "01001000",
    4206 => "01001000",
    4207 => "01001000",
    4208 => "01001000",
    4209 => "01001000",
    4210 => "01001000",
    4211 => "01001000",
    4212 => "01001000",
    4213 => "01001000",
    4214 => "01001000",
    4215 => "01001000",
    4216 => "01001000",
    4217 => "01001000",
    4218 => "01001000",
    4219 => "01001000",
    4220 => "01001000",
    4221 => "01001000",
    4222 => "01001000",
    4223 => "01001000",
    4224 => "01001000",
    4225 => "01001000",
    4226 => "01001000",
    4227 => "01001000",
    4228 => "01001000",
    4229 => "01001000",
    4230 => "01001000",
    4231 => "01001000",
    4232 => "01000111",
    4233 => "01000111",
    4234 => "01000111",
    4235 => "01000111",
    4236 => "01000111",
    4237 => "01000111",
    4238 => "01000111",
    4239 => "01000111",
    4240 => "01000111",
    4241 => "01000111",
    4242 => "01000111",
    4243 => "01000111",
    4244 => "01000111",
    4245 => "01000111",
    4246 => "01000111",
    4247 => "01000111",
    4248 => "01000111",
    4249 => "01000111",
    4250 => "01000111",
    4251 => "01000111",
    4252 => "01000111",
    4253 => "01000111",
    4254 => "01000111",
    4255 => "01000111",
    4256 => "01000111",
    4257 => "01000111",
    4258 => "01000111",
    4259 => "01000111",
    4260 => "01000111",
    4261 => "01000111",
    4262 => "01000111",
    4263 => "01000111",
    4264 => "01000111",
    4265 => "01000111",
    4266 => "01000111",
    4267 => "01000111",
    4268 => "01000111",
    4269 => "01000111",
    4270 => "01000111",
    4271 => "01000111",
    4272 => "01000111",
    4273 => "01000111",
    4274 => "01000111",
    4275 => "01000111",
    4276 => "01000111",
    4277 => "01000111",
    4278 => "01000111",
    4279 => "01000110",
    4280 => "01000110",
    4281 => "01000110",
    4282 => "01000110",
    4283 => "01000110",
    4284 => "01000110",
    4285 => "01000110",
    4286 => "01000110",
    4287 => "01000110",
    4288 => "01000110",
    4289 => "01000110",
    4290 => "01000110",
    4291 => "01000110",
    4292 => "01000110",
    4293 => "01000110",
    4294 => "01000110",
    4295 => "01000110",
    4296 => "01000110",
    4297 => "01000110",
    4298 => "01000110",
    4299 => "01000110",
    4300 => "01000110",
    4301 => "01000110",
    4302 => "01000110",
    4303 => "01000110",
    4304 => "01000110",
    4305 => "01000110",
    4306 => "01000110",
    4307 => "01000110",
    4308 => "01000110",
    4309 => "01000110",
    4310 => "01000110",
    4311 => "01000110",
    4312 => "01000110",
    4313 => "01000110",
    4314 => "01000110",
    4315 => "01000110",
    4316 => "01000110",
    4317 => "01000110",
    4318 => "01000110",
    4319 => "01000110",
    4320 => "01000110",
    4321 => "01000110",
    4322 => "01000110",
    4323 => "01000110",
    4324 => "01000110",
    4325 => "01000101",
    4326 => "01000101",
    4327 => "01000101",
    4328 => "01000101",
    4329 => "01000101",
    4330 => "01000101",
    4331 => "01000101",
    4332 => "01000101",
    4333 => "01000101",
    4334 => "01000101",
    4335 => "01000101",
    4336 => "01000101",
    4337 => "01000101",
    4338 => "01000101",
    4339 => "01000101",
    4340 => "01000101",
    4341 => "01000101",
    4342 => "01000101",
    4343 => "01000101",
    4344 => "01000101",
    4345 => "01000101",
    4346 => "01000101",
    4347 => "01000101",
    4348 => "01000101",
    4349 => "01000101",
    4350 => "01000101",
    4351 => "01000101",
    4352 => "01000101",
    4353 => "01000101",
    4354 => "01000101",
    4355 => "01000101",
    4356 => "01000101",
    4357 => "01000101",
    4358 => "01000101",
    4359 => "01000101",
    4360 => "01000101",
    4361 => "01000101",
    4362 => "01000101",
    4363 => "01000101",
    4364 => "01000101",
    4365 => "01000101",
    4366 => "01000101",
    4367 => "01000101",
    4368 => "01000101",
    4369 => "01000101",
    4370 => "01000101",
    4371 => "01000101",
    4372 => "01000100",
    4373 => "01000100",
    4374 => "01000100",
    4375 => "01000100",
    4376 => "01000100",
    4377 => "01000100",
    4378 => "01000100",
    4379 => "01000100",
    4380 => "01000100",
    4381 => "01000100",
    4382 => "01000100",
    4383 => "01000100",
    4384 => "01000100",
    4385 => "01000100",
    4386 => "01000100",
    4387 => "01000100",
    4388 => "01000100",
    4389 => "01000100",
    4390 => "01000100",
    4391 => "01000100",
    4392 => "01000100",
    4393 => "01000100",
    4394 => "01000100",
    4395 => "01000100",
    4396 => "01000100",
    4397 => "01000100",
    4398 => "01000100",
    4399 => "01000100",
    4400 => "01000100",
    4401 => "01000100",
    4402 => "01000100",
    4403 => "01000100",
    4404 => "01000100",
    4405 => "01000100",
    4406 => "01000100",
    4407 => "01000100",
    4408 => "01000100",
    4409 => "01000100",
    4410 => "01000100",
    4411 => "01000100",
    4412 => "01000100",
    4413 => "01000100",
    4414 => "01000100",
    4415 => "01000100",
    4416 => "01000100",
    4417 => "01000100",
    4418 => "01000011",
    4419 => "01000011",
    4420 => "01000011",
    4421 => "01000011",
    4422 => "01000011",
    4423 => "01000011",
    4424 => "01000011",
    4425 => "01000011",
    4426 => "01000011",
    4427 => "01000011",
    4428 => "01000011",
    4429 => "01000011",
    4430 => "01000011",
    4431 => "01000011",
    4432 => "01000011",
    4433 => "01000011",
    4434 => "01000011",
    4435 => "01000011",
    4436 => "01000011",
    4437 => "01000011",
    4438 => "01000011",
    4439 => "01000011",
    4440 => "01000011",
    4441 => "01000011",
    4442 => "01000011",
    4443 => "01000011",
    4444 => "01000011",
    4445 => "01000011",
    4446 => "01000011",
    4447 => "01000011",
    4448 => "01000011",
    4449 => "01000011",
    4450 => "01000011",
    4451 => "01000011",
    4452 => "01000011",
    4453 => "01000011",
    4454 => "01000011",
    4455 => "01000011",
    4456 => "01000011",
    4457 => "01000011",
    4458 => "01000011",
    4459 => "01000011",
    4460 => "01000011",
    4461 => "01000011",
    4462 => "01000011",
    4463 => "01000011",
    4464 => "01000011",
    4465 => "01000011",
    4466 => "01000010",
    4467 => "01000010",
    4468 => "01000010",
    4469 => "01000010",
    4470 => "01000010",
    4471 => "01000010",
    4472 => "01000010",
    4473 => "01000010",
    4474 => "01000010",
    4475 => "01000010",
    4476 => "01000010",
    4477 => "01000010",
    4478 => "01000010",
    4479 => "01000010",
    4480 => "01000010",
    4481 => "01000010",
    4482 => "01000010",
    4483 => "01000010",
    4484 => "01000010",
    4485 => "01000010",
    4486 => "01000010",
    4487 => "01000010",
    4488 => "01000010",
    4489 => "01000010",
    4490 => "01000010",
    4491 => "01000010",
    4492 => "01000010",
    4493 => "01000010",
    4494 => "01000010",
    4495 => "01000010",
    4496 => "01000010",
    4497 => "01000010",
    4498 => "01000010",
    4499 => "01000010",
    4500 => "01000010",
    4501 => "01000010",
    4502 => "01000010",
    4503 => "01000010",
    4504 => "01000010",
    4505 => "01000010",
    4506 => "01000010",
    4507 => "01000010",
    4508 => "01000010",
    4509 => "01000010",
    4510 => "01000010",
    4511 => "01000010",
    4512 => "01000010",
    4513 => "01000001",
    4514 => "01000001",
    4515 => "01000001",
    4516 => "01000001",
    4517 => "01000001",
    4518 => "01000001",
    4519 => "01000001",
    4520 => "01000001",
    4521 => "01000001",
    4522 => "01000001",
    4523 => "01000001",
    4524 => "01000001",
    4525 => "01000001",
    4526 => "01000001",
    4527 => "01000001",
    4528 => "01000001",
    4529 => "01000001",
    4530 => "01000001",
    4531 => "01000001",
    4532 => "01000001",
    4533 => "01000001",
    4534 => "01000001",
    4535 => "01000001",
    4536 => "01000001",
    4537 => "01000001",
    4538 => "01000001",
    4539 => "01000001",
    4540 => "01000001",
    4541 => "01000001",
    4542 => "01000001",
    4543 => "01000001",
    4544 => "01000001",
    4545 => "01000001",
    4546 => "01000001",
    4547 => "01000001",
    4548 => "01000001",
    4549 => "01000001",
    4550 => "01000001",
    4551 => "01000001",
    4552 => "01000001",
    4553 => "01000001",
    4554 => "01000001",
    4555 => "01000001",
    4556 => "01000001",
    4557 => "01000001",
    4558 => "01000001",
    4559 => "01000001",
    4560 => "01000001",
    4561 => "01000000",
    4562 => "01000000",
    4563 => "01000000",
    4564 => "01000000",
    4565 => "01000000",
    4566 => "01000000",
    4567 => "01000000",
    4568 => "01000000",
    4569 => "01000000",
    4570 => "01000000",
    4571 => "01000000",
    4572 => "01000000",
    4573 => "01000000",
    4574 => "01000000",
    4575 => "01000000",
    4576 => "01000000",
    4577 => "01000000",
    4578 => "01000000",
    4579 => "01000000",
    4580 => "01000000",
    4581 => "01000000",
    4582 => "01000000",
    4583 => "01000000",
    4584 => "01000000",
    4585 => "01000000",
    4586 => "01000000",
    4587 => "01000000",
    4588 => "01000000",
    4589 => "01000000",
    4590 => "01000000",
    4591 => "01000000",
    4592 => "01000000",
    4593 => "01000000",
    4594 => "01000000",
    4595 => "01000000",
    4596 => "01000000",
    4597 => "01000000",
    4598 => "01000000",
    4599 => "01000000",
    4600 => "01000000",
    4601 => "01000000",
    4602 => "01000000",
    4603 => "01000000",
    4604 => "01000000",
    4605 => "01000000",
    4606 => "01000000",
    4607 => "01000000",
    4608 => "00111111",
    4609 => "00111111",
    4610 => "00111111",
    4611 => "00111111",
    4612 => "00111111",
    4613 => "00111111",
    4614 => "00111111",
    4615 => "00111111",
    4616 => "00111111",
    4617 => "00111111",
    4618 => "00111111",
    4619 => "00111111",
    4620 => "00111111",
    4621 => "00111111",
    4622 => "00111111",
    4623 => "00111111",
    4624 => "00111111",
    4625 => "00111111",
    4626 => "00111111",
    4627 => "00111111",
    4628 => "00111111",
    4629 => "00111111",
    4630 => "00111111",
    4631 => "00111111",
    4632 => "00111111",
    4633 => "00111111",
    4634 => "00111111",
    4635 => "00111111",
    4636 => "00111111",
    4637 => "00111111",
    4638 => "00111111",
    4639 => "00111111",
    4640 => "00111111",
    4641 => "00111111",
    4642 => "00111111",
    4643 => "00111111",
    4644 => "00111111",
    4645 => "00111111",
    4646 => "00111111",
    4647 => "00111111",
    4648 => "00111111",
    4649 => "00111111",
    4650 => "00111111",
    4651 => "00111111",
    4652 => "00111111",
    4653 => "00111111",
    4654 => "00111111",
    4655 => "00111111",
    4656 => "00111111",
    4657 => "00111110",
    4658 => "00111110",
    4659 => "00111110",
    4660 => "00111110",
    4661 => "00111110",
    4662 => "00111110",
    4663 => "00111110",
    4664 => "00111110",
    4665 => "00111110",
    4666 => "00111110",
    4667 => "00111110",
    4668 => "00111110",
    4669 => "00111110",
    4670 => "00111110",
    4671 => "00111110",
    4672 => "00111110",
    4673 => "00111110",
    4674 => "00111110",
    4675 => "00111110",
    4676 => "00111110",
    4677 => "00111110",
    4678 => "00111110",
    4679 => "00111110",
    4680 => "00111110",
    4681 => "00111110",
    4682 => "00111110",
    4683 => "00111110",
    4684 => "00111110",
    4685 => "00111110",
    4686 => "00111110",
    4687 => "00111110",
    4688 => "00111110",
    4689 => "00111110",
    4690 => "00111110",
    4691 => "00111110",
    4692 => "00111110",
    4693 => "00111110",
    4694 => "00111110",
    4695 => "00111110",
    4696 => "00111110",
    4697 => "00111110",
    4698 => "00111110",
    4699 => "00111110",
    4700 => "00111110",
    4701 => "00111110",
    4702 => "00111110",
    4703 => "00111110",
    4704 => "00111110",
    4705 => "00111101",
    4706 => "00111101",
    4707 => "00111101",
    4708 => "00111101",
    4709 => "00111101",
    4710 => "00111101",
    4711 => "00111101",
    4712 => "00111101",
    4713 => "00111101",
    4714 => "00111101",
    4715 => "00111101",
    4716 => "00111101",
    4717 => "00111101",
    4718 => "00111101",
    4719 => "00111101",
    4720 => "00111101",
    4721 => "00111101",
    4722 => "00111101",
    4723 => "00111101",
    4724 => "00111101",
    4725 => "00111101",
    4726 => "00111101",
    4727 => "00111101",
    4728 => "00111101",
    4729 => "00111101",
    4730 => "00111101",
    4731 => "00111101",
    4732 => "00111101",
    4733 => "00111101",
    4734 => "00111101",
    4735 => "00111101",
    4736 => "00111101",
    4737 => "00111101",
    4738 => "00111101",
    4739 => "00111101",
    4740 => "00111101",
    4741 => "00111101",
    4742 => "00111101",
    4743 => "00111101",
    4744 => "00111101",
    4745 => "00111101",
    4746 => "00111101",
    4747 => "00111101",
    4748 => "00111101",
    4749 => "00111101",
    4750 => "00111101",
    4751 => "00111101",
    4752 => "00111101",
    4753 => "00111101",
    4754 => "00111100",
    4755 => "00111100",
    4756 => "00111100",
    4757 => "00111100",
    4758 => "00111100",
    4759 => "00111100",
    4760 => "00111100",
    4761 => "00111100",
    4762 => "00111100",
    4763 => "00111100",
    4764 => "00111100",
    4765 => "00111100",
    4766 => "00111100",
    4767 => "00111100",
    4768 => "00111100",
    4769 => "00111100",
    4770 => "00111100",
    4771 => "00111100",
    4772 => "00111100",
    4773 => "00111100",
    4774 => "00111100",
    4775 => "00111100",
    4776 => "00111100",
    4777 => "00111100",
    4778 => "00111100",
    4779 => "00111100",
    4780 => "00111100",
    4781 => "00111100",
    4782 => "00111100",
    4783 => "00111100",
    4784 => "00111100",
    4785 => "00111100",
    4786 => "00111100",
    4787 => "00111100",
    4788 => "00111100",
    4789 => "00111100",
    4790 => "00111100",
    4791 => "00111100",
    4792 => "00111100",
    4793 => "00111100",
    4794 => "00111100",
    4795 => "00111100",
    4796 => "00111100",
    4797 => "00111100",
    4798 => "00111100",
    4799 => "00111100",
    4800 => "00111100",
    4801 => "00111100",
    4802 => "00111011",
    4803 => "00111011",
    4804 => "00111011",
    4805 => "00111011",
    4806 => "00111011",
    4807 => "00111011",
    4808 => "00111011",
    4809 => "00111011",
    4810 => "00111011",
    4811 => "00111011",
    4812 => "00111011",
    4813 => "00111011",
    4814 => "00111011",
    4815 => "00111011",
    4816 => "00111011",
    4817 => "00111011",
    4818 => "00111011",
    4819 => "00111011",
    4820 => "00111011",
    4821 => "00111011",
    4822 => "00111011",
    4823 => "00111011",
    4824 => "00111011",
    4825 => "00111011",
    4826 => "00111011",
    4827 => "00111011",
    4828 => "00111011",
    4829 => "00111011",
    4830 => "00111011",
    4831 => "00111011",
    4832 => "00111011",
    4833 => "00111011",
    4834 => "00111011",
    4835 => "00111011",
    4836 => "00111011",
    4837 => "00111011",
    4838 => "00111011",
    4839 => "00111011",
    4840 => "00111011",
    4841 => "00111011",
    4842 => "00111011",
    4843 => "00111011",
    4844 => "00111011",
    4845 => "00111011",
    4846 => "00111011",
    4847 => "00111011",
    4848 => "00111011",
    4849 => "00111011",
    4850 => "00111011",
    4851 => "00111011",
    4852 => "00111010",
    4853 => "00111010",
    4854 => "00111010",
    4855 => "00111010",
    4856 => "00111010",
    4857 => "00111010",
    4858 => "00111010",
    4859 => "00111010",
    4860 => "00111010",
    4861 => "00111010",
    4862 => "00111010",
    4863 => "00111010",
    4864 => "00111010",
    4865 => "00111010",
    4866 => "00111010",
    4867 => "00111010",
    4868 => "00111010",
    4869 => "00111010",
    4870 => "00111010",
    4871 => "00111010",
    4872 => "00111010",
    4873 => "00111010",
    4874 => "00111010",
    4875 => "00111010",
    4876 => "00111010",
    4877 => "00111010",
    4878 => "00111010",
    4879 => "00111010",
    4880 => "00111010",
    4881 => "00111010",
    4882 => "00111010",
    4883 => "00111010",
    4884 => "00111010",
    4885 => "00111010",
    4886 => "00111010",
    4887 => "00111010",
    4888 => "00111010",
    4889 => "00111010",
    4890 => "00111010",
    4891 => "00111010",
    4892 => "00111010",
    4893 => "00111010",
    4894 => "00111010",
    4895 => "00111010",
    4896 => "00111010",
    4897 => "00111010",
    4898 => "00111010",
    4899 => "00111010",
    4900 => "00111010",
    4901 => "00111001",
    4902 => "00111001",
    4903 => "00111001",
    4904 => "00111001",
    4905 => "00111001",
    4906 => "00111001",
    4907 => "00111001",
    4908 => "00111001",
    4909 => "00111001",
    4910 => "00111001",
    4911 => "00111001",
    4912 => "00111001",
    4913 => "00111001",
    4914 => "00111001",
    4915 => "00111001",
    4916 => "00111001",
    4917 => "00111001",
    4918 => "00111001",
    4919 => "00111001",
    4920 => "00111001",
    4921 => "00111001",
    4922 => "00111001",
    4923 => "00111001",
    4924 => "00111001",
    4925 => "00111001",
    4926 => "00111001",
    4927 => "00111001",
    4928 => "00111001",
    4929 => "00111001",
    4930 => "00111001",
    4931 => "00111001",
    4932 => "00111001",
    4933 => "00111001",
    4934 => "00111001",
    4935 => "00111001",
    4936 => "00111001",
    4937 => "00111001",
    4938 => "00111001",
    4939 => "00111001",
    4940 => "00111001",
    4941 => "00111001",
    4942 => "00111001",
    4943 => "00111001",
    4944 => "00111001",
    4945 => "00111001",
    4946 => "00111001",
    4947 => "00111001",
    4948 => "00111001",
    4949 => "00111001",
    4950 => "00111001",
    4951 => "00111000",
    4952 => "00111000",
    4953 => "00111000",
    4954 => "00111000",
    4955 => "00111000",
    4956 => "00111000",
    4957 => "00111000",
    4958 => "00111000",
    4959 => "00111000",
    4960 => "00111000",
    4961 => "00111000",
    4962 => "00111000",
    4963 => "00111000",
    4964 => "00111000",
    4965 => "00111000",
    4966 => "00111000",
    4967 => "00111000",
    4968 => "00111000",
    4969 => "00111000",
    4970 => "00111000",
    4971 => "00111000",
    4972 => "00111000",
    4973 => "00111000",
    4974 => "00111000",
    4975 => "00111000",
    4976 => "00111000",
    4977 => "00111000",
    4978 => "00111000",
    4979 => "00111000",
    4980 => "00111000",
    4981 => "00111000",
    4982 => "00111000",
    4983 => "00111000",
    4984 => "00111000",
    4985 => "00111000",
    4986 => "00111000",
    4987 => "00111000",
    4988 => "00111000",
    4989 => "00111000",
    4990 => "00111000",
    4991 => "00111000",
    4992 => "00111000",
    4993 => "00111000",
    4994 => "00111000",
    4995 => "00111000",
    4996 => "00111000",
    4997 => "00111000",
    4998 => "00111000",
    4999 => "00111000",
    5000 => "00110111",
    5001 => "00110111",
    5002 => "00110111",
    5003 => "00110111",
    5004 => "00110111",
    5005 => "00110111",
    5006 => "00110111",
    5007 => "00110111",
    5008 => "00110111",
    5009 => "00110111",
    5010 => "00110111",
    5011 => "00110111",
    5012 => "00110111",
    5013 => "00110111",
    5014 => "00110111",
    5015 => "00110111",
    5016 => "00110111",
    5017 => "00110111",
    5018 => "00110111",
    5019 => "00110111",
    5020 => "00110111",
    5021 => "00110111",
    5022 => "00110111",
    5023 => "00110111",
    5024 => "00110111",
    5025 => "00110111",
    5026 => "00110111",
    5027 => "00110111",
    5028 => "00110111",
    5029 => "00110111",
    5030 => "00110111",
    5031 => "00110111",
    5032 => "00110111",
    5033 => "00110111",
    5034 => "00110111",
    5035 => "00110111",
    5036 => "00110111",
    5037 => "00110111",
    5038 => "00110111",
    5039 => "00110111",
    5040 => "00110111",
    5041 => "00110111",
    5042 => "00110111",
    5043 => "00110111",
    5044 => "00110111",
    5045 => "00110111",
    5046 => "00110111",
    5047 => "00110111",
    5048 => "00110111",
    5049 => "00110111",
    5050 => "00110111",
    5051 => "00110110",
    5052 => "00110110",
    5053 => "00110110",
    5054 => "00110110",
    5055 => "00110110",
    5056 => "00110110",
    5057 => "00110110",
    5058 => "00110110",
    5059 => "00110110",
    5060 => "00110110",
    5061 => "00110110",
    5062 => "00110110",
    5063 => "00110110",
    5064 => "00110110",
    5065 => "00110110",
    5066 => "00110110",
    5067 => "00110110",
    5068 => "00110110",
    5069 => "00110110",
    5070 => "00110110",
    5071 => "00110110",
    5072 => "00110110",
    5073 => "00110110",
    5074 => "00110110",
    5075 => "00110110",
    5076 => "00110110",
    5077 => "00110110",
    5078 => "00110110",
    5079 => "00110110",
    5080 => "00110110",
    5081 => "00110110",
    5082 => "00110110",
    5083 => "00110110",
    5084 => "00110110",
    5085 => "00110110",
    5086 => "00110110",
    5087 => "00110110",
    5088 => "00110110",
    5089 => "00110110",
    5090 => "00110110",
    5091 => "00110110",
    5092 => "00110110",
    5093 => "00110110",
    5094 => "00110110",
    5095 => "00110110",
    5096 => "00110110",
    5097 => "00110110",
    5098 => "00110110",
    5099 => "00110110",
    5100 => "00110110",
    5101 => "00110101",
    5102 => "00110101",
    5103 => "00110101",
    5104 => "00110101",
    5105 => "00110101",
    5106 => "00110101",
    5107 => "00110101",
    5108 => "00110101",
    5109 => "00110101",
    5110 => "00110101",
    5111 => "00110101",
    5112 => "00110101",
    5113 => "00110101",
    5114 => "00110101",
    5115 => "00110101",
    5116 => "00110101",
    5117 => "00110101",
    5118 => "00110101",
    5119 => "00110101",
    5120 => "00110101",
    5121 => "00110101",
    5122 => "00110101",
    5123 => "00110101",
    5124 => "00110101",
    5125 => "00110101",
    5126 => "00110101",
    5127 => "00110101",
    5128 => "00110101",
    5129 => "00110101",
    5130 => "00110101",
    5131 => "00110101",
    5132 => "00110101",
    5133 => "00110101",
    5134 => "00110101",
    5135 => "00110101",
    5136 => "00110101",
    5137 => "00110101",
    5138 => "00110101",
    5139 => "00110101",
    5140 => "00110101",
    5141 => "00110101",
    5142 => "00110101",
    5143 => "00110101",
    5144 => "00110101",
    5145 => "00110101",
    5146 => "00110101",
    5147 => "00110101",
    5148 => "00110101",
    5149 => "00110101",
    5150 => "00110101",
    5151 => "00110101",
    5152 => "00110100",
    5153 => "00110100",
    5154 => "00110100",
    5155 => "00110100",
    5156 => "00110100",
    5157 => "00110100",
    5158 => "00110100",
    5159 => "00110100",
    5160 => "00110100",
    5161 => "00110100",
    5162 => "00110100",
    5163 => "00110100",
    5164 => "00110100",
    5165 => "00110100",
    5166 => "00110100",
    5167 => "00110100",
    5168 => "00110100",
    5169 => "00110100",
    5170 => "00110100",
    5171 => "00110100",
    5172 => "00110100",
    5173 => "00110100",
    5174 => "00110100",
    5175 => "00110100",
    5176 => "00110100",
    5177 => "00110100",
    5178 => "00110100",
    5179 => "00110100",
    5180 => "00110100",
    5181 => "00110100",
    5182 => "00110100",
    5183 => "00110100",
    5184 => "00110100",
    5185 => "00110100",
    5186 => "00110100",
    5187 => "00110100",
    5188 => "00110100",
    5189 => "00110100",
    5190 => "00110100",
    5191 => "00110100",
    5192 => "00110100",
    5193 => "00110100",
    5194 => "00110100",
    5195 => "00110100",
    5196 => "00110100",
    5197 => "00110100",
    5198 => "00110100",
    5199 => "00110100",
    5200 => "00110100",
    5201 => "00110100",
    5202 => "00110011",
    5203 => "00110011",
    5204 => "00110011",
    5205 => "00110011",
    5206 => "00110011",
    5207 => "00110011",
    5208 => "00110011",
    5209 => "00110011",
    5210 => "00110011",
    5211 => "00110011",
    5212 => "00110011",
    5213 => "00110011",
    5214 => "00110011",
    5215 => "00110011",
    5216 => "00110011",
    5217 => "00110011",
    5218 => "00110011",
    5219 => "00110011",
    5220 => "00110011",
    5221 => "00110011",
    5222 => "00110011",
    5223 => "00110011",
    5224 => "00110011",
    5225 => "00110011",
    5226 => "00110011",
    5227 => "00110011",
    5228 => "00110011",
    5229 => "00110011",
    5230 => "00110011",
    5231 => "00110011",
    5232 => "00110011",
    5233 => "00110011",
    5234 => "00110011",
    5235 => "00110011",
    5236 => "00110011",
    5237 => "00110011",
    5238 => "00110011",
    5239 => "00110011",
    5240 => "00110011",
    5241 => "00110011",
    5242 => "00110011",
    5243 => "00110011",
    5244 => "00110011",
    5245 => "00110011",
    5246 => "00110011",
    5247 => "00110011",
    5248 => "00110011",
    5249 => "00110011",
    5250 => "00110011",
    5251 => "00110011",
    5252 => "00110011",
    5253 => "00110011",
    5254 => "00110010",
    5255 => "00110010",
    5256 => "00110010",
    5257 => "00110010",
    5258 => "00110010",
    5259 => "00110010",
    5260 => "00110010",
    5261 => "00110010",
    5262 => "00110010",
    5263 => "00110010",
    5264 => "00110010",
    5265 => "00110010",
    5266 => "00110010",
    5267 => "00110010",
    5268 => "00110010",
    5269 => "00110010",
    5270 => "00110010",
    5271 => "00110010",
    5272 => "00110010",
    5273 => "00110010",
    5274 => "00110010",
    5275 => "00110010",
    5276 => "00110010",
    5277 => "00110010",
    5278 => "00110010",
    5279 => "00110010",
    5280 => "00110010",
    5281 => "00110010",
    5282 => "00110010",
    5283 => "00110010",
    5284 => "00110010",
    5285 => "00110010",
    5286 => "00110010",
    5287 => "00110010",
    5288 => "00110010",
    5289 => "00110010",
    5290 => "00110010",
    5291 => "00110010",
    5292 => "00110010",
    5293 => "00110010",
    5294 => "00110010",
    5295 => "00110010",
    5296 => "00110010",
    5297 => "00110010",
    5298 => "00110010",
    5299 => "00110010",
    5300 => "00110010",
    5301 => "00110010",
    5302 => "00110010",
    5303 => "00110010",
    5304 => "00110010",
    5305 => "00110001",
    5306 => "00110001",
    5307 => "00110001",
    5308 => "00110001",
    5309 => "00110001",
    5310 => "00110001",
    5311 => "00110001",
    5312 => "00110001",
    5313 => "00110001",
    5314 => "00110001",
    5315 => "00110001",
    5316 => "00110001",
    5317 => "00110001",
    5318 => "00110001",
    5319 => "00110001",
    5320 => "00110001",
    5321 => "00110001",
    5322 => "00110001",
    5323 => "00110001",
    5324 => "00110001",
    5325 => "00110001",
    5326 => "00110001",
    5327 => "00110001",
    5328 => "00110001",
    5329 => "00110001",
    5330 => "00110001",
    5331 => "00110001",
    5332 => "00110001",
    5333 => "00110001",
    5334 => "00110001",
    5335 => "00110001",
    5336 => "00110001",
    5337 => "00110001",
    5338 => "00110001",
    5339 => "00110001",
    5340 => "00110001",
    5341 => "00110001",
    5342 => "00110001",
    5343 => "00110001",
    5344 => "00110001",
    5345 => "00110001",
    5346 => "00110001",
    5347 => "00110001",
    5348 => "00110001",
    5349 => "00110001",
    5350 => "00110001",
    5351 => "00110001",
    5352 => "00110001",
    5353 => "00110001",
    5354 => "00110001",
    5355 => "00110001",
    5356 => "00110001",
    5357 => "00110000",
    5358 => "00110000",
    5359 => "00110000",
    5360 => "00110000",
    5361 => "00110000",
    5362 => "00110000",
    5363 => "00110000",
    5364 => "00110000",
    5365 => "00110000",
    5366 => "00110000",
    5367 => "00110000",
    5368 => "00110000",
    5369 => "00110000",
    5370 => "00110000",
    5371 => "00110000",
    5372 => "00110000",
    5373 => "00110000",
    5374 => "00110000",
    5375 => "00110000",
    5376 => "00110000",
    5377 => "00110000",
    5378 => "00110000",
    5379 => "00110000",
    5380 => "00110000",
    5381 => "00110000",
    5382 => "00110000",
    5383 => "00110000",
    5384 => "00110000",
    5385 => "00110000",
    5386 => "00110000",
    5387 => "00110000",
    5388 => "00110000",
    5389 => "00110000",
    5390 => "00110000",
    5391 => "00110000",
    5392 => "00110000",
    5393 => "00110000",
    5394 => "00110000",
    5395 => "00110000",
    5396 => "00110000",
    5397 => "00110000",
    5398 => "00110000",
    5399 => "00110000",
    5400 => "00110000",
    5401 => "00110000",
    5402 => "00110000",
    5403 => "00110000",
    5404 => "00110000",
    5405 => "00110000",
    5406 => "00110000",
    5407 => "00110000",
    5408 => "00101111",
    5409 => "00101111",
    5410 => "00101111",
    5411 => "00101111",
    5412 => "00101111",
    5413 => "00101111",
    5414 => "00101111",
    5415 => "00101111",
    5416 => "00101111",
    5417 => "00101111",
    5418 => "00101111",
    5419 => "00101111",
    5420 => "00101111",
    5421 => "00101111",
    5422 => "00101111",
    5423 => "00101111",
    5424 => "00101111",
    5425 => "00101111",
    5426 => "00101111",
    5427 => "00101111",
    5428 => "00101111",
    5429 => "00101111",
    5430 => "00101111",
    5431 => "00101111",
    5432 => "00101111",
    5433 => "00101111",
    5434 => "00101111",
    5435 => "00101111",
    5436 => "00101111",
    5437 => "00101111",
    5438 => "00101111",
    5439 => "00101111",
    5440 => "00101111",
    5441 => "00101111",
    5442 => "00101111",
    5443 => "00101111",
    5444 => "00101111",
    5445 => "00101111",
    5446 => "00101111",
    5447 => "00101111",
    5448 => "00101111",
    5449 => "00101111",
    5450 => "00101111",
    5451 => "00101111",
    5452 => "00101111",
    5453 => "00101111",
    5454 => "00101111",
    5455 => "00101111",
    5456 => "00101111",
    5457 => "00101111",
    5458 => "00101111",
    5459 => "00101111",
    5460 => "00101111",
    5461 => "00101110",
    5462 => "00101110",
    5463 => "00101110",
    5464 => "00101110",
    5465 => "00101110",
    5466 => "00101110",
    5467 => "00101110",
    5468 => "00101110",
    5469 => "00101110",
    5470 => "00101110",
    5471 => "00101110",
    5472 => "00101110",
    5473 => "00101110",
    5474 => "00101110",
    5475 => "00101110",
    5476 => "00101110",
    5477 => "00101110",
    5478 => "00101110",
    5479 => "00101110",
    5480 => "00101110",
    5481 => "00101110",
    5482 => "00101110",
    5483 => "00101110",
    5484 => "00101110",
    5485 => "00101110",
    5486 => "00101110",
    5487 => "00101110",
    5488 => "00101110",
    5489 => "00101110",
    5490 => "00101110",
    5491 => "00101110",
    5492 => "00101110",
    5493 => "00101110",
    5494 => "00101110",
    5495 => "00101110",
    5496 => "00101110",
    5497 => "00101110",
    5498 => "00101110",
    5499 => "00101110",
    5500 => "00101110",
    5501 => "00101110",
    5502 => "00101110",
    5503 => "00101110",
    5504 => "00101110",
    5505 => "00101110",
    5506 => "00101110",
    5507 => "00101110",
    5508 => "00101110",
    5509 => "00101110",
    5510 => "00101110",
    5511 => "00101110",
    5512 => "00101110",
    5513 => "00101101",
    5514 => "00101101",
    5515 => "00101101",
    5516 => "00101101",
    5517 => "00101101",
    5518 => "00101101",
    5519 => "00101101",
    5520 => "00101101",
    5521 => "00101101",
    5522 => "00101101",
    5523 => "00101101",
    5524 => "00101101",
    5525 => "00101101",
    5526 => "00101101",
    5527 => "00101101",
    5528 => "00101101",
    5529 => "00101101",
    5530 => "00101101",
    5531 => "00101101",
    5532 => "00101101",
    5533 => "00101101",
    5534 => "00101101",
    5535 => "00101101",
    5536 => "00101101",
    5537 => "00101101",
    5538 => "00101101",
    5539 => "00101101",
    5540 => "00101101",
    5541 => "00101101",
    5542 => "00101101",
    5543 => "00101101",
    5544 => "00101101",
    5545 => "00101101",
    5546 => "00101101",
    5547 => "00101101",
    5548 => "00101101",
    5549 => "00101101",
    5550 => "00101101",
    5551 => "00101101",
    5552 => "00101101",
    5553 => "00101101",
    5554 => "00101101",
    5555 => "00101101",
    5556 => "00101101",
    5557 => "00101101",
    5558 => "00101101",
    5559 => "00101101",
    5560 => "00101101",
    5561 => "00101101",
    5562 => "00101101",
    5563 => "00101101",
    5564 => "00101101",
    5565 => "00101101",
    5566 => "00101100",
    5567 => "00101100",
    5568 => "00101100",
    5569 => "00101100",
    5570 => "00101100",
    5571 => "00101100",
    5572 => "00101100",
    5573 => "00101100",
    5574 => "00101100",
    5575 => "00101100",
    5576 => "00101100",
    5577 => "00101100",
    5578 => "00101100",
    5579 => "00101100",
    5580 => "00101100",
    5581 => "00101100",
    5582 => "00101100",
    5583 => "00101100",
    5584 => "00101100",
    5585 => "00101100",
    5586 => "00101100",
    5587 => "00101100",
    5588 => "00101100",
    5589 => "00101100",
    5590 => "00101100",
    5591 => "00101100",
    5592 => "00101100",
    5593 => "00101100",
    5594 => "00101100",
    5595 => "00101100",
    5596 => "00101100",
    5597 => "00101100",
    5598 => "00101100",
    5599 => "00101100",
    5600 => "00101100",
    5601 => "00101100",
    5602 => "00101100",
    5603 => "00101100",
    5604 => "00101100",
    5605 => "00101100",
    5606 => "00101100",
    5607 => "00101100",
    5608 => "00101100",
    5609 => "00101100",
    5610 => "00101100",
    5611 => "00101100",
    5612 => "00101100",
    5613 => "00101100",
    5614 => "00101100",
    5615 => "00101100",
    5616 => "00101100",
    5617 => "00101100",
    5618 => "00101011",
    5619 => "00101011",
    5620 => "00101011",
    5621 => "00101011",
    5622 => "00101011",
    5623 => "00101011",
    5624 => "00101011",
    5625 => "00101011",
    5626 => "00101011",
    5627 => "00101011",
    5628 => "00101011",
    5629 => "00101011",
    5630 => "00101011",
    5631 => "00101011",
    5632 => "00101011",
    5633 => "00101011",
    5634 => "00101011",
    5635 => "00101011",
    5636 => "00101011",
    5637 => "00101011",
    5638 => "00101011",
    5639 => "00101011",
    5640 => "00101011",
    5641 => "00101011",
    5642 => "00101011",
    5643 => "00101011",
    5644 => "00101011",
    5645 => "00101011",
    5646 => "00101011",
    5647 => "00101011",
    5648 => "00101011",
    5649 => "00101011",
    5650 => "00101011",
    5651 => "00101011",
    5652 => "00101011",
    5653 => "00101011",
    5654 => "00101011",
    5655 => "00101011",
    5656 => "00101011",
    5657 => "00101011",
    5658 => "00101011",
    5659 => "00101011",
    5660 => "00101011",
    5661 => "00101011",
    5662 => "00101011",
    5663 => "00101011",
    5664 => "00101011",
    5665 => "00101011",
    5666 => "00101011",
    5667 => "00101011",
    5668 => "00101011",
    5669 => "00101011",
    5670 => "00101011",
    5671 => "00101011",
    5672 => "00101010",
    5673 => "00101010",
    5674 => "00101010",
    5675 => "00101010",
    5676 => "00101010",
    5677 => "00101010",
    5678 => "00101010",
    5679 => "00101010",
    5680 => "00101010",
    5681 => "00101010",
    5682 => "00101010",
    5683 => "00101010",
    5684 => "00101010",
    5685 => "00101010",
    5686 => "00101010",
    5687 => "00101010",
    5688 => "00101010",
    5689 => "00101010",
    5690 => "00101010",
    5691 => "00101010",
    5692 => "00101010",
    5693 => "00101010",
    5694 => "00101010",
    5695 => "00101010",
    5696 => "00101010",
    5697 => "00101010",
    5698 => "00101010",
    5699 => "00101010",
    5700 => "00101010",
    5701 => "00101010",
    5702 => "00101010",
    5703 => "00101010",
    5704 => "00101010",
    5705 => "00101010",
    5706 => "00101010",
    5707 => "00101010",
    5708 => "00101010",
    5709 => "00101010",
    5710 => "00101010",
    5711 => "00101010",
    5712 => "00101010",
    5713 => "00101010",
    5714 => "00101010",
    5715 => "00101010",
    5716 => "00101010",
    5717 => "00101010",
    5718 => "00101010",
    5719 => "00101010",
    5720 => "00101010",
    5721 => "00101010",
    5722 => "00101010",
    5723 => "00101010",
    5724 => "00101010",
    5725 => "00101001",
    5726 => "00101001",
    5727 => "00101001",
    5728 => "00101001",
    5729 => "00101001",
    5730 => "00101001",
    5731 => "00101001",
    5732 => "00101001",
    5733 => "00101001",
    5734 => "00101001",
    5735 => "00101001",
    5736 => "00101001",
    5737 => "00101001",
    5738 => "00101001",
    5739 => "00101001",
    5740 => "00101001",
    5741 => "00101001",
    5742 => "00101001",
    5743 => "00101001",
    5744 => "00101001",
    5745 => "00101001",
    5746 => "00101001",
    5747 => "00101001",
    5748 => "00101001",
    5749 => "00101001",
    5750 => "00101001",
    5751 => "00101001",
    5752 => "00101001",
    5753 => "00101001",
    5754 => "00101001",
    5755 => "00101001",
    5756 => "00101001",
    5757 => "00101001",
    5758 => "00101001",
    5759 => "00101001",
    5760 => "00101001",
    5761 => "00101001",
    5762 => "00101001",
    5763 => "00101001",
    5764 => "00101001",
    5765 => "00101001",
    5766 => "00101001",
    5767 => "00101001",
    5768 => "00101001",
    5769 => "00101001",
    5770 => "00101001",
    5771 => "00101001",
    5772 => "00101001",
    5773 => "00101001",
    5774 => "00101001",
    5775 => "00101001",
    5776 => "00101001",
    5777 => "00101001",
    5778 => "00101001",
    5779 => "00101000",
    5780 => "00101000",
    5781 => "00101000",
    5782 => "00101000",
    5783 => "00101000",
    5784 => "00101000",
    5785 => "00101000",
    5786 => "00101000",
    5787 => "00101000",
    5788 => "00101000",
    5789 => "00101000",
    5790 => "00101000",
    5791 => "00101000",
    5792 => "00101000",
    5793 => "00101000",
    5794 => "00101000",
    5795 => "00101000",
    5796 => "00101000",
    5797 => "00101000",
    5798 => "00101000",
    5799 => "00101000",
    5800 => "00101000",
    5801 => "00101000",
    5802 => "00101000",
    5803 => "00101000",
    5804 => "00101000",
    5805 => "00101000",
    5806 => "00101000",
    5807 => "00101000",
    5808 => "00101000",
    5809 => "00101000",
    5810 => "00101000",
    5811 => "00101000",
    5812 => "00101000",
    5813 => "00101000",
    5814 => "00101000",
    5815 => "00101000",
    5816 => "00101000",
    5817 => "00101000",
    5818 => "00101000",
    5819 => "00101000",
    5820 => "00101000",
    5821 => "00101000",
    5822 => "00101000",
    5823 => "00101000",
    5824 => "00101000",
    5825 => "00101000",
    5826 => "00101000",
    5827 => "00101000",
    5828 => "00101000",
    5829 => "00101000",
    5830 => "00101000",
    5831 => "00101000",
    5832 => "00100111",
    5833 => "00100111",
    5834 => "00100111",
    5835 => "00100111",
    5836 => "00100111",
    5837 => "00100111",
    5838 => "00100111",
    5839 => "00100111",
    5840 => "00100111",
    5841 => "00100111",
    5842 => "00100111",
    5843 => "00100111",
    5844 => "00100111",
    5845 => "00100111",
    5846 => "00100111",
    5847 => "00100111",
    5848 => "00100111",
    5849 => "00100111",
    5850 => "00100111",
    5851 => "00100111",
    5852 => "00100111",
    5853 => "00100111",
    5854 => "00100111",
    5855 => "00100111",
    5856 => "00100111",
    5857 => "00100111",
    5858 => "00100111",
    5859 => "00100111",
    5860 => "00100111",
    5861 => "00100111",
    5862 => "00100111",
    5863 => "00100111",
    5864 => "00100111",
    5865 => "00100111",
    5866 => "00100111",
    5867 => "00100111",
    5868 => "00100111",
    5869 => "00100111",
    5870 => "00100111",
    5871 => "00100111",
    5872 => "00100111",
    5873 => "00100111",
    5874 => "00100111",
    5875 => "00100111",
    5876 => "00100111",
    5877 => "00100111",
    5878 => "00100111",
    5879 => "00100111",
    5880 => "00100111",
    5881 => "00100111",
    5882 => "00100111",
    5883 => "00100111",
    5884 => "00100111",
    5885 => "00100111",
    5886 => "00100111",
    5887 => "00100110",
    5888 => "00100110",
    5889 => "00100110",
    5890 => "00100110",
    5891 => "00100110",
    5892 => "00100110",
    5893 => "00100110",
    5894 => "00100110",
    5895 => "00100110",
    5896 => "00100110",
    5897 => "00100110",
    5898 => "00100110",
    5899 => "00100110",
    5900 => "00100110",
    5901 => "00100110",
    5902 => "00100110",
    5903 => "00100110",
    5904 => "00100110",
    5905 => "00100110",
    5906 => "00100110",
    5907 => "00100110",
    5908 => "00100110",
    5909 => "00100110",
    5910 => "00100110",
    5911 => "00100110",
    5912 => "00100110",
    5913 => "00100110",
    5914 => "00100110",
    5915 => "00100110",
    5916 => "00100110",
    5917 => "00100110",
    5918 => "00100110",
    5919 => "00100110",
    5920 => "00100110",
    5921 => "00100110",
    5922 => "00100110",
    5923 => "00100110",
    5924 => "00100110",
    5925 => "00100110",
    5926 => "00100110",
    5927 => "00100110",
    5928 => "00100110",
    5929 => "00100110",
    5930 => "00100110",
    5931 => "00100110",
    5932 => "00100110",
    5933 => "00100110",
    5934 => "00100110",
    5935 => "00100110",
    5936 => "00100110",
    5937 => "00100110",
    5938 => "00100110",
    5939 => "00100110",
    5940 => "00100110",
    5941 => "00100101",
    5942 => "00100101",
    5943 => "00100101",
    5944 => "00100101",
    5945 => "00100101",
    5946 => "00100101",
    5947 => "00100101",
    5948 => "00100101",
    5949 => "00100101",
    5950 => "00100101",
    5951 => "00100101",
    5952 => "00100101",
    5953 => "00100101",
    5954 => "00100101",
    5955 => "00100101",
    5956 => "00100101",
    5957 => "00100101",
    5958 => "00100101",
    5959 => "00100101",
    5960 => "00100101",
    5961 => "00100101",
    5962 => "00100101",
    5963 => "00100101",
    5964 => "00100101",
    5965 => "00100101",
    5966 => "00100101",
    5967 => "00100101",
    5968 => "00100101",
    5969 => "00100101",
    5970 => "00100101",
    5971 => "00100101",
    5972 => "00100101",
    5973 => "00100101",
    5974 => "00100101",
    5975 => "00100101",
    5976 => "00100101",
    5977 => "00100101",
    5978 => "00100101",
    5979 => "00100101",
    5980 => "00100101",
    5981 => "00100101",
    5982 => "00100101",
    5983 => "00100101",
    5984 => "00100101",
    5985 => "00100101",
    5986 => "00100101",
    5987 => "00100101",
    5988 => "00100101",
    5989 => "00100101",
    5990 => "00100101",
    5991 => "00100101",
    5992 => "00100101",
    5993 => "00100101",
    5994 => "00100101",
    5995 => "00100101",
    5996 => "00100100",
    5997 => "00100100",
    5998 => "00100100",
    5999 => "00100100",
    6000 => "00100100",
    6001 => "00100100",
    6002 => "00100100",
    6003 => "00100100",
    6004 => "00100100",
    6005 => "00100100",
    6006 => "00100100",
    6007 => "00100100",
    6008 => "00100100",
    6009 => "00100100",
    6010 => "00100100",
    6011 => "00100100",
    6012 => "00100100",
    6013 => "00100100",
    6014 => "00100100",
    6015 => "00100100",
    6016 => "00100100",
    6017 => "00100100",
    6018 => "00100100",
    6019 => "00100100",
    6020 => "00100100",
    6021 => "00100100",
    6022 => "00100100",
    6023 => "00100100",
    6024 => "00100100",
    6025 => "00100100",
    6026 => "00100100",
    6027 => "00100100",
    6028 => "00100100",
    6029 => "00100100",
    6030 => "00100100",
    6031 => "00100100",
    6032 => "00100100",
    6033 => "00100100",
    6034 => "00100100",
    6035 => "00100100",
    6036 => "00100100",
    6037 => "00100100",
    6038 => "00100100",
    6039 => "00100100",
    6040 => "00100100",
    6041 => "00100100",
    6042 => "00100100",
    6043 => "00100100",
    6044 => "00100100",
    6045 => "00100100",
    6046 => "00100100",
    6047 => "00100100",
    6048 => "00100100",
    6049 => "00100100",
    6050 => "00100011",
    6051 => "00100011",
    6052 => "00100011",
    6053 => "00100011",
    6054 => "00100011",
    6055 => "00100011",
    6056 => "00100011",
    6057 => "00100011",
    6058 => "00100011",
    6059 => "00100011",
    6060 => "00100011",
    6061 => "00100011",
    6062 => "00100011",
    6063 => "00100011",
    6064 => "00100011",
    6065 => "00100011",
    6066 => "00100011",
    6067 => "00100011",
    6068 => "00100011",
    6069 => "00100011",
    6070 => "00100011",
    6071 => "00100011",
    6072 => "00100011",
    6073 => "00100011",
    6074 => "00100011",
    6075 => "00100011",
    6076 => "00100011",
    6077 => "00100011",
    6078 => "00100011",
    6079 => "00100011",
    6080 => "00100011",
    6081 => "00100011",
    6082 => "00100011",
    6083 => "00100011",
    6084 => "00100011",
    6085 => "00100011",
    6086 => "00100011",
    6087 => "00100011",
    6088 => "00100011",
    6089 => "00100011",
    6090 => "00100011",
    6091 => "00100011",
    6092 => "00100011",
    6093 => "00100011",
    6094 => "00100011",
    6095 => "00100011",
    6096 => "00100011",
    6097 => "00100011",
    6098 => "00100011",
    6099 => "00100011",
    6100 => "00100011",
    6101 => "00100011",
    6102 => "00100011",
    6103 => "00100011",
    6104 => "00100011",
    6105 => "00100011",
    6106 => "00100010",
    6107 => "00100010",
    6108 => "00100010",
    6109 => "00100010",
    6110 => "00100010",
    6111 => "00100010",
    6112 => "00100010",
    6113 => "00100010",
    6114 => "00100010",
    6115 => "00100010",
    6116 => "00100010",
    6117 => "00100010",
    6118 => "00100010",
    6119 => "00100010",
    6120 => "00100010",
    6121 => "00100010",
    6122 => "00100010",
    6123 => "00100010",
    6124 => "00100010",
    6125 => "00100010",
    6126 => "00100010",
    6127 => "00100010",
    6128 => "00100010",
    6129 => "00100010",
    6130 => "00100010",
    6131 => "00100010",
    6132 => "00100010",
    6133 => "00100010",
    6134 => "00100010",
    6135 => "00100010",
    6136 => "00100010",
    6137 => "00100010",
    6138 => "00100010",
    6139 => "00100010",
    6140 => "00100010",
    6141 => "00100010",
    6142 => "00100010",
    6143 => "00100010",
    6144 => "00100010",
    6145 => "00100010",
    6146 => "00100010",
    6147 => "00100010",
    6148 => "00100010",
    6149 => "00100010",
    6150 => "00100010",
    6151 => "00100010",
    6152 => "00100010",
    6153 => "00100010",
    6154 => "00100010",
    6155 => "00100010",
    6156 => "00100010",
    6157 => "00100010",
    6158 => "00100010",
    6159 => "00100010",
    6160 => "00100010",
    6161 => "00100001",
    6162 => "00100001",
    6163 => "00100001",
    6164 => "00100001",
    6165 => "00100001",
    6166 => "00100001",
    6167 => "00100001",
    6168 => "00100001",
    6169 => "00100001",
    6170 => "00100001",
    6171 => "00100001",
    6172 => "00100001",
    6173 => "00100001",
    6174 => "00100001",
    6175 => "00100001",
    6176 => "00100001",
    6177 => "00100001",
    6178 => "00100001",
    6179 => "00100001",
    6180 => "00100001",
    6181 => "00100001",
    6182 => "00100001",
    6183 => "00100001",
    6184 => "00100001",
    6185 => "00100001",
    6186 => "00100001",
    6187 => "00100001",
    6188 => "00100001",
    6189 => "00100001",
    6190 => "00100001",
    6191 => "00100001",
    6192 => "00100001",
    6193 => "00100001",
    6194 => "00100001",
    6195 => "00100001",
    6196 => "00100001",
    6197 => "00100001",
    6198 => "00100001",
    6199 => "00100001",
    6200 => "00100001",
    6201 => "00100001",
    6202 => "00100001",
    6203 => "00100001",
    6204 => "00100001",
    6205 => "00100001",
    6206 => "00100001",
    6207 => "00100001",
    6208 => "00100001",
    6209 => "00100001",
    6210 => "00100001",
    6211 => "00100001",
    6212 => "00100001",
    6213 => "00100001",
    6214 => "00100001",
    6215 => "00100001",
    6216 => "00100001",
    6217 => "00100000",
    6218 => "00100000",
    6219 => "00100000",
    6220 => "00100000",
    6221 => "00100000",
    6222 => "00100000",
    6223 => "00100000",
    6224 => "00100000",
    6225 => "00100000",
    6226 => "00100000",
    6227 => "00100000",
    6228 => "00100000",
    6229 => "00100000",
    6230 => "00100000",
    6231 => "00100000",
    6232 => "00100000",
    6233 => "00100000",
    6234 => "00100000",
    6235 => "00100000",
    6236 => "00100000",
    6237 => "00100000",
    6238 => "00100000",
    6239 => "00100000",
    6240 => "00100000",
    6241 => "00100000",
    6242 => "00100000",
    6243 => "00100000",
    6244 => "00100000",
    6245 => "00100000",
    6246 => "00100000",
    6247 => "00100000",
    6248 => "00100000",
    6249 => "00100000",
    6250 => "00100000",
    6251 => "00100000",
    6252 => "00100000",
    6253 => "00100000",
    6254 => "00100000",
    6255 => "00100000",
    6256 => "00100000",
    6257 => "00100000",
    6258 => "00100000",
    6259 => "00100000",
    6260 => "00100000",
    6261 => "00100000",
    6262 => "00100000",
    6263 => "00100000",
    6264 => "00100000",
    6265 => "00100000",
    6266 => "00100000",
    6267 => "00100000",
    6268 => "00100000",
    6269 => "00100000",
    6270 => "00100000",
    6271 => "00100000",
    6272 => "00011111",
    6273 => "00011111",
    6274 => "00011111",
    6275 => "00011111",
    6276 => "00011111",
    6277 => "00011111",
    6278 => "00011111",
    6279 => "00011111",
    6280 => "00011111",
    6281 => "00011111",
    6282 => "00011111",
    6283 => "00011111",
    6284 => "00011111",
    6285 => "00011111",
    6286 => "00011111",
    6287 => "00011111",
    6288 => "00011111",
    6289 => "00011111",
    6290 => "00011111",
    6291 => "00011111",
    6292 => "00011111",
    6293 => "00011111",
    6294 => "00011111",
    6295 => "00011111",
    6296 => "00011111",
    6297 => "00011111",
    6298 => "00011111",
    6299 => "00011111",
    6300 => "00011111",
    6301 => "00011111",
    6302 => "00011111",
    6303 => "00011111",
    6304 => "00011111",
    6305 => "00011111",
    6306 => "00011111",
    6307 => "00011111",
    6308 => "00011111",
    6309 => "00011111",
    6310 => "00011111",
    6311 => "00011111",
    6312 => "00011111",
    6313 => "00011111",
    6314 => "00011111",
    6315 => "00011111",
    6316 => "00011111",
    6317 => "00011111",
    6318 => "00011111",
    6319 => "00011111",
    6320 => "00011111",
    6321 => "00011111",
    6322 => "00011111",
    6323 => "00011111",
    6324 => "00011111",
    6325 => "00011111",
    6326 => "00011111",
    6327 => "00011111",
    6328 => "00011111",
    6329 => "00011110",
    6330 => "00011110",
    6331 => "00011110",
    6332 => "00011110",
    6333 => "00011110",
    6334 => "00011110",
    6335 => "00011110",
    6336 => "00011110",
    6337 => "00011110",
    6338 => "00011110",
    6339 => "00011110",
    6340 => "00011110",
    6341 => "00011110",
    6342 => "00011110",
    6343 => "00011110",
    6344 => "00011110",
    6345 => "00011110",
    6346 => "00011110",
    6347 => "00011110",
    6348 => "00011110",
    6349 => "00011110",
    6350 => "00011110",
    6351 => "00011110",
    6352 => "00011110",
    6353 => "00011110",
    6354 => "00011110",
    6355 => "00011110",
    6356 => "00011110",
    6357 => "00011110",
    6358 => "00011110",
    6359 => "00011110",
    6360 => "00011110",
    6361 => "00011110",
    6362 => "00011110",
    6363 => "00011110",
    6364 => "00011110",
    6365 => "00011110",
    6366 => "00011110",
    6367 => "00011110",
    6368 => "00011110",
    6369 => "00011110",
    6370 => "00011110",
    6371 => "00011110",
    6372 => "00011110",
    6373 => "00011110",
    6374 => "00011110",
    6375 => "00011110",
    6376 => "00011110",
    6377 => "00011110",
    6378 => "00011110",
    6379 => "00011110",
    6380 => "00011110",
    6381 => "00011110",
    6382 => "00011110",
    6383 => "00011110",
    6384 => "00011110",
    6385 => "00011101",
    6386 => "00011101",
    6387 => "00011101",
    6388 => "00011101",
    6389 => "00011101",
    6390 => "00011101",
    6391 => "00011101",
    6392 => "00011101",
    6393 => "00011101",
    6394 => "00011101",
    6395 => "00011101",
    6396 => "00011101",
    6397 => "00011101",
    6398 => "00011101",
    6399 => "00011101",
    6400 => "00011101",
    6401 => "00011101",
    6402 => "00011101",
    6403 => "00011101",
    6404 => "00011101",
    6405 => "00011101",
    6406 => "00011101",
    6407 => "00011101",
    6408 => "00011101",
    6409 => "00011101",
    6410 => "00011101",
    6411 => "00011101",
    6412 => "00011101",
    6413 => "00011101",
    6414 => "00011101",
    6415 => "00011101",
    6416 => "00011101",
    6417 => "00011101",
    6418 => "00011101",
    6419 => "00011101",
    6420 => "00011101",
    6421 => "00011101",
    6422 => "00011101",
    6423 => "00011101",
    6424 => "00011101",
    6425 => "00011101",
    6426 => "00011101",
    6427 => "00011101",
    6428 => "00011101",
    6429 => "00011101",
    6430 => "00011101",
    6431 => "00011101",
    6432 => "00011101",
    6433 => "00011101",
    6434 => "00011101",
    6435 => "00011101",
    6436 => "00011101",
    6437 => "00011101",
    6438 => "00011101",
    6439 => "00011101",
    6440 => "00011101",
    6441 => "00011101",
    6442 => "00011100",
    6443 => "00011100",
    6444 => "00011100",
    6445 => "00011100",
    6446 => "00011100",
    6447 => "00011100",
    6448 => "00011100",
    6449 => "00011100",
    6450 => "00011100",
    6451 => "00011100",
    6452 => "00011100",
    6453 => "00011100",
    6454 => "00011100",
    6455 => "00011100",
    6456 => "00011100",
    6457 => "00011100",
    6458 => "00011100",
    6459 => "00011100",
    6460 => "00011100",
    6461 => "00011100",
    6462 => "00011100",
    6463 => "00011100",
    6464 => "00011100",
    6465 => "00011100",
    6466 => "00011100",
    6467 => "00011100",
    6468 => "00011100",
    6469 => "00011100",
    6470 => "00011100",
    6471 => "00011100",
    6472 => "00011100",
    6473 => "00011100",
    6474 => "00011100",
    6475 => "00011100",
    6476 => "00011100",
    6477 => "00011100",
    6478 => "00011100",
    6479 => "00011100",
    6480 => "00011100",
    6481 => "00011100",
    6482 => "00011100",
    6483 => "00011100",
    6484 => "00011100",
    6485 => "00011100",
    6486 => "00011100",
    6487 => "00011100",
    6488 => "00011100",
    6489 => "00011100",
    6490 => "00011100",
    6491 => "00011100",
    6492 => "00011100",
    6493 => "00011100",
    6494 => "00011100",
    6495 => "00011100",
    6496 => "00011100",
    6497 => "00011100",
    6498 => "00011011",
    6499 => "00011011",
    6500 => "00011011",
    6501 => "00011011",
    6502 => "00011011",
    6503 => "00011011",
    6504 => "00011011",
    6505 => "00011011",
    6506 => "00011011",
    6507 => "00011011",
    6508 => "00011011",
    6509 => "00011011",
    6510 => "00011011",
    6511 => "00011011",
    6512 => "00011011",
    6513 => "00011011",
    6514 => "00011011",
    6515 => "00011011",
    6516 => "00011011",
    6517 => "00011011",
    6518 => "00011011",
    6519 => "00011011",
    6520 => "00011011",
    6521 => "00011011",
    6522 => "00011011",
    6523 => "00011011",
    6524 => "00011011",
    6525 => "00011011",
    6526 => "00011011",
    6527 => "00011011",
    6528 => "00011011",
    6529 => "00011011",
    6530 => "00011011",
    6531 => "00011011",
    6532 => "00011011",
    6533 => "00011011",
    6534 => "00011011",
    6535 => "00011011",
    6536 => "00011011",
    6537 => "00011011",
    6538 => "00011011",
    6539 => "00011011",
    6540 => "00011011",
    6541 => "00011011",
    6542 => "00011011",
    6543 => "00011011",
    6544 => "00011011",
    6545 => "00011011",
    6546 => "00011011",
    6547 => "00011011",
    6548 => "00011011",
    6549 => "00011011",
    6550 => "00011011",
    6551 => "00011011",
    6552 => "00011011",
    6553 => "00011011",
    6554 => "00011011",
    6555 => "00011011",
    6556 => "00011010",
    6557 => "00011010",
    6558 => "00011010",
    6559 => "00011010",
    6560 => "00011010",
    6561 => "00011010",
    6562 => "00011010",
    6563 => "00011010",
    6564 => "00011010",
    6565 => "00011010",
    6566 => "00011010",
    6567 => "00011010",
    6568 => "00011010",
    6569 => "00011010",
    6570 => "00011010",
    6571 => "00011010",
    6572 => "00011010",
    6573 => "00011010",
    6574 => "00011010",
    6575 => "00011010",
    6576 => "00011010",
    6577 => "00011010",
    6578 => "00011010",
    6579 => "00011010",
    6580 => "00011010",
    6581 => "00011010",
    6582 => "00011010",
    6583 => "00011010",
    6584 => "00011010",
    6585 => "00011010",
    6586 => "00011010",
    6587 => "00011010",
    6588 => "00011010",
    6589 => "00011010",
    6590 => "00011010",
    6591 => "00011010",
    6592 => "00011010",
    6593 => "00011010",
    6594 => "00011010",
    6595 => "00011010",
    6596 => "00011010",
    6597 => "00011010",
    6598 => "00011010",
    6599 => "00011010",
    6600 => "00011010",
    6601 => "00011010",
    6602 => "00011010",
    6603 => "00011010",
    6604 => "00011010",
    6605 => "00011010",
    6606 => "00011010",
    6607 => "00011010",
    6608 => "00011010",
    6609 => "00011010",
    6610 => "00011010",
    6611 => "00011010",
    6612 => "00011010",
    6613 => "00011001",
    6614 => "00011001",
    6615 => "00011001",
    6616 => "00011001",
    6617 => "00011001",
    6618 => "00011001",
    6619 => "00011001",
    6620 => "00011001",
    6621 => "00011001",
    6622 => "00011001",
    6623 => "00011001",
    6624 => "00011001",
    6625 => "00011001",
    6626 => "00011001",
    6627 => "00011001",
    6628 => "00011001",
    6629 => "00011001",
    6630 => "00011001",
    6631 => "00011001",
    6632 => "00011001",
    6633 => "00011001",
    6634 => "00011001",
    6635 => "00011001",
    6636 => "00011001",
    6637 => "00011001",
    6638 => "00011001",
    6639 => "00011001",
    6640 => "00011001",
    6641 => "00011001",
    6642 => "00011001",
    6643 => "00011001",
    6644 => "00011001",
    6645 => "00011001",
    6646 => "00011001",
    6647 => "00011001",
    6648 => "00011001",
    6649 => "00011001",
    6650 => "00011001",
    6651 => "00011001",
    6652 => "00011001",
    6653 => "00011001",
    6654 => "00011001",
    6655 => "00011001",
    6656 => "00011001",
    6657 => "00011001",
    6658 => "00011001",
    6659 => "00011001",
    6660 => "00011001",
    6661 => "00011001",
    6662 => "00011001",
    6663 => "00011001",
    6664 => "00011001",
    6665 => "00011001",
    6666 => "00011001",
    6667 => "00011001",
    6668 => "00011001",
    6669 => "00011001",
    6670 => "00011001",
    6671 => "00011000",
    6672 => "00011000",
    6673 => "00011000",
    6674 => "00011000",
    6675 => "00011000",
    6676 => "00011000",
    6677 => "00011000",
    6678 => "00011000",
    6679 => "00011000",
    6680 => "00011000",
    6681 => "00011000",
    6682 => "00011000",
    6683 => "00011000",
    6684 => "00011000",
    6685 => "00011000",
    6686 => "00011000",
    6687 => "00011000",
    6688 => "00011000",
    6689 => "00011000",
    6690 => "00011000",
    6691 => "00011000",
    6692 => "00011000",
    6693 => "00011000",
    6694 => "00011000",
    6695 => "00011000",
    6696 => "00011000",
    6697 => "00011000",
    6698 => "00011000",
    6699 => "00011000",
    6700 => "00011000",
    6701 => "00011000",
    6702 => "00011000",
    6703 => "00011000",
    6704 => "00011000",
    6705 => "00011000",
    6706 => "00011000",
    6707 => "00011000",
    6708 => "00011000",
    6709 => "00011000",
    6710 => "00011000",
    6711 => "00011000",
    6712 => "00011000",
    6713 => "00011000",
    6714 => "00011000",
    6715 => "00011000",
    6716 => "00011000",
    6717 => "00011000",
    6718 => "00011000",
    6719 => "00011000",
    6720 => "00011000",
    6721 => "00011000",
    6722 => "00011000",
    6723 => "00011000",
    6724 => "00011000",
    6725 => "00011000",
    6726 => "00011000",
    6727 => "00011000",
    6728 => "00010111",
    6729 => "00010111",
    6730 => "00010111",
    6731 => "00010111",
    6732 => "00010111",
    6733 => "00010111",
    6734 => "00010111",
    6735 => "00010111",
    6736 => "00010111",
    6737 => "00010111",
    6738 => "00010111",
    6739 => "00010111",
    6740 => "00010111",
    6741 => "00010111",
    6742 => "00010111",
    6743 => "00010111",
    6744 => "00010111",
    6745 => "00010111",
    6746 => "00010111",
    6747 => "00010111",
    6748 => "00010111",
    6749 => "00010111",
    6750 => "00010111",
    6751 => "00010111",
    6752 => "00010111",
    6753 => "00010111",
    6754 => "00010111",
    6755 => "00010111",
    6756 => "00010111",
    6757 => "00010111",
    6758 => "00010111",
    6759 => "00010111",
    6760 => "00010111",
    6761 => "00010111",
    6762 => "00010111",
    6763 => "00010111",
    6764 => "00010111",
    6765 => "00010111",
    6766 => "00010111",
    6767 => "00010111",
    6768 => "00010111",
    6769 => "00010111",
    6770 => "00010111",
    6771 => "00010111",
    6772 => "00010111",
    6773 => "00010111",
    6774 => "00010111",
    6775 => "00010111",
    6776 => "00010111",
    6777 => "00010111",
    6778 => "00010111",
    6779 => "00010111",
    6780 => "00010111",
    6781 => "00010111",
    6782 => "00010111",
    6783 => "00010111",
    6784 => "00010111",
    6785 => "00010111",
    6786 => "00010111",
    6787 => "00010110",
    6788 => "00010110",
    6789 => "00010110",
    6790 => "00010110",
    6791 => "00010110",
    6792 => "00010110",
    6793 => "00010110",
    6794 => "00010110",
    6795 => "00010110",
    6796 => "00010110",
    6797 => "00010110",
    6798 => "00010110",
    6799 => "00010110",
    6800 => "00010110",
    6801 => "00010110",
    6802 => "00010110",
    6803 => "00010110",
    6804 => "00010110",
    6805 => "00010110",
    6806 => "00010110",
    6807 => "00010110",
    6808 => "00010110",
    6809 => "00010110",
    6810 => "00010110",
    6811 => "00010110",
    6812 => "00010110",
    6813 => "00010110",
    6814 => "00010110",
    6815 => "00010110",
    6816 => "00010110",
    6817 => "00010110",
    6818 => "00010110",
    6819 => "00010110",
    6820 => "00010110",
    6821 => "00010110",
    6822 => "00010110",
    6823 => "00010110",
    6824 => "00010110",
    6825 => "00010110",
    6826 => "00010110",
    6827 => "00010110",
    6828 => "00010110",
    6829 => "00010110",
    6830 => "00010110",
    6831 => "00010110",
    6832 => "00010110",
    6833 => "00010110",
    6834 => "00010110",
    6835 => "00010110",
    6836 => "00010110",
    6837 => "00010110",
    6838 => "00010110",
    6839 => "00010110",
    6840 => "00010110",
    6841 => "00010110",
    6842 => "00010110",
    6843 => "00010110",
    6844 => "00010110",
    6845 => "00010101",
    6846 => "00010101",
    6847 => "00010101",
    6848 => "00010101",
    6849 => "00010101",
    6850 => "00010101",
    6851 => "00010101",
    6852 => "00010101",
    6853 => "00010101",
    6854 => "00010101",
    6855 => "00010101",
    6856 => "00010101",
    6857 => "00010101",
    6858 => "00010101",
    6859 => "00010101",
    6860 => "00010101",
    6861 => "00010101",
    6862 => "00010101",
    6863 => "00010101",
    6864 => "00010101",
    6865 => "00010101",
    6866 => "00010101",
    6867 => "00010101",
    6868 => "00010101",
    6869 => "00010101",
    6870 => "00010101",
    6871 => "00010101",
    6872 => "00010101",
    6873 => "00010101",
    6874 => "00010101",
    6875 => "00010101",
    6876 => "00010101",
    6877 => "00010101",
    6878 => "00010101",
    6879 => "00010101",
    6880 => "00010101",
    6881 => "00010101",
    6882 => "00010101",
    6883 => "00010101",
    6884 => "00010101",
    6885 => "00010101",
    6886 => "00010101",
    6887 => "00010101",
    6888 => "00010101",
    6889 => "00010101",
    6890 => "00010101",
    6891 => "00010101",
    6892 => "00010101",
    6893 => "00010101",
    6894 => "00010101",
    6895 => "00010101",
    6896 => "00010101",
    6897 => "00010101",
    6898 => "00010101",
    6899 => "00010101",
    6900 => "00010101",
    6901 => "00010101",
    6902 => "00010101",
    6903 => "00010101",
    6904 => "00010100",
    6905 => "00010100",
    6906 => "00010100",
    6907 => "00010100",
    6908 => "00010100",
    6909 => "00010100",
    6910 => "00010100",
    6911 => "00010100",
    6912 => "00010100",
    6913 => "00010100",
    6914 => "00010100",
    6915 => "00010100",
    6916 => "00010100",
    6917 => "00010100",
    6918 => "00010100",
    6919 => "00010100",
    6920 => "00010100",
    6921 => "00010100",
    6922 => "00010100",
    6923 => "00010100",
    6924 => "00010100",
    6925 => "00010100",
    6926 => "00010100",
    6927 => "00010100",
    6928 => "00010100",
    6929 => "00010100",
    6930 => "00010100",
    6931 => "00010100",
    6932 => "00010100",
    6933 => "00010100",
    6934 => "00010100",
    6935 => "00010100",
    6936 => "00010100",
    6937 => "00010100",
    6938 => "00010100",
    6939 => "00010100",
    6940 => "00010100",
    6941 => "00010100",
    6942 => "00010100",
    6943 => "00010100",
    6944 => "00010100",
    6945 => "00010100",
    6946 => "00010100",
    6947 => "00010100",
    6948 => "00010100",
    6949 => "00010100",
    6950 => "00010100",
    6951 => "00010100",
    6952 => "00010100",
    6953 => "00010100",
    6954 => "00010100",
    6955 => "00010100",
    6956 => "00010100",
    6957 => "00010100",
    6958 => "00010100",
    6959 => "00010100",
    6960 => "00010100",
    6961 => "00010100",
    6962 => "00010011",
    6963 => "00010011",
    6964 => "00010011",
    6965 => "00010011",
    6966 => "00010011",
    6967 => "00010011",
    6968 => "00010011",
    6969 => "00010011",
    6970 => "00010011",
    6971 => "00010011",
    6972 => "00010011",
    6973 => "00010011",
    6974 => "00010011",
    6975 => "00010011",
    6976 => "00010011",
    6977 => "00010011",
    6978 => "00010011",
    6979 => "00010011",
    6980 => "00010011",
    6981 => "00010011",
    6982 => "00010011",
    6983 => "00010011",
    6984 => "00010011",
    6985 => "00010011",
    6986 => "00010011",
    6987 => "00010011",
    6988 => "00010011",
    6989 => "00010011",
    6990 => "00010011",
    6991 => "00010011",
    6992 => "00010011",
    6993 => "00010011",
    6994 => "00010011",
    6995 => "00010011",
    6996 => "00010011",
    6997 => "00010011",
    6998 => "00010011",
    6999 => "00010011",
    7000 => "00010011",
    7001 => "00010011",
    7002 => "00010011",
    7003 => "00010011",
    7004 => "00010011",
    7005 => "00010011",
    7006 => "00010011",
    7007 => "00010011",
    7008 => "00010011",
    7009 => "00010011",
    7010 => "00010011",
    7011 => "00010011",
    7012 => "00010011",
    7013 => "00010011",
    7014 => "00010011",
    7015 => "00010011",
    7016 => "00010011",
    7017 => "00010011",
    7018 => "00010011",
    7019 => "00010011",
    7020 => "00010011",
    7021 => "00010011",
    7022 => "00010010",
    7023 => "00010010",
    7024 => "00010010",
    7025 => "00010010",
    7026 => "00010010",
    7027 => "00010010",
    7028 => "00010010",
    7029 => "00010010",
    7030 => "00010010",
    7031 => "00010010",
    7032 => "00010010",
    7033 => "00010010",
    7034 => "00010010",
    7035 => "00010010",
    7036 => "00010010",
    7037 => "00010010",
    7038 => "00010010",
    7039 => "00010010",
    7040 => "00010010",
    7041 => "00010010",
    7042 => "00010010",
    7043 => "00010010",
    7044 => "00010010",
    7045 => "00010010",
    7046 => "00010010",
    7047 => "00010010",
    7048 => "00010010",
    7049 => "00010010",
    7050 => "00010010",
    7051 => "00010010",
    7052 => "00010010",
    7053 => "00010010",
    7054 => "00010010",
    7055 => "00010010",
    7056 => "00010010",
    7057 => "00010010",
    7058 => "00010010",
    7059 => "00010010",
    7060 => "00010010",
    7061 => "00010010",
    7062 => "00010010",
    7063 => "00010010",
    7064 => "00010010",
    7065 => "00010010",
    7066 => "00010010",
    7067 => "00010010",
    7068 => "00010010",
    7069 => "00010010",
    7070 => "00010010",
    7071 => "00010010",
    7072 => "00010010",
    7073 => "00010010",
    7074 => "00010010",
    7075 => "00010010",
    7076 => "00010010",
    7077 => "00010010",
    7078 => "00010010",
    7079 => "00010010",
    7080 => "00010010",
    7081 => "00010001",
    7082 => "00010001",
    7083 => "00010001",
    7084 => "00010001",
    7085 => "00010001",
    7086 => "00010001",
    7087 => "00010001",
    7088 => "00010001",
    7089 => "00010001",
    7090 => "00010001",
    7091 => "00010001",
    7092 => "00010001",
    7093 => "00010001",
    7094 => "00010001",
    7095 => "00010001",
    7096 => "00010001",
    7097 => "00010001",
    7098 => "00010001",
    7099 => "00010001",
    7100 => "00010001",
    7101 => "00010001",
    7102 => "00010001",
    7103 => "00010001",
    7104 => "00010001",
    7105 => "00010001",
    7106 => "00010001",
    7107 => "00010001",
    7108 => "00010001",
    7109 => "00010001",
    7110 => "00010001",
    7111 => "00010001",
    7112 => "00010001",
    7113 => "00010001",
    7114 => "00010001",
    7115 => "00010001",
    7116 => "00010001",
    7117 => "00010001",
    7118 => "00010001",
    7119 => "00010001",
    7120 => "00010001",
    7121 => "00010001",
    7122 => "00010001",
    7123 => "00010001",
    7124 => "00010001",
    7125 => "00010001",
    7126 => "00010001",
    7127 => "00010001",
    7128 => "00010001",
    7129 => "00010001",
    7130 => "00010001",
    7131 => "00010001",
    7132 => "00010001",
    7133 => "00010001",
    7134 => "00010001",
    7135 => "00010001",
    7136 => "00010001",
    7137 => "00010001",
    7138 => "00010001",
    7139 => "00010001",
    7140 => "00010001",
    7141 => "00010000",
    7142 => "00010000",
    7143 => "00010000",
    7144 => "00010000",
    7145 => "00010000",
    7146 => "00010000",
    7147 => "00010000",
    7148 => "00010000",
    7149 => "00010000",
    7150 => "00010000",
    7151 => "00010000",
    7152 => "00010000",
    7153 => "00010000",
    7154 => "00010000",
    7155 => "00010000",
    7156 => "00010000",
    7157 => "00010000",
    7158 => "00010000",
    7159 => "00010000",
    7160 => "00010000",
    7161 => "00010000",
    7162 => "00010000",
    7163 => "00010000",
    7164 => "00010000",
    7165 => "00010000",
    7166 => "00010000",
    7167 => "00010000",
    7168 => "00010000",
    7169 => "00010000",
    7170 => "00010000",
    7171 => "00010000",
    7172 => "00010000",
    7173 => "00010000",
    7174 => "00010000",
    7175 => "00010000",
    7176 => "00010000",
    7177 => "00010000",
    7178 => "00010000",
    7179 => "00010000",
    7180 => "00010000",
    7181 => "00010000",
    7182 => "00010000",
    7183 => "00010000",
    7184 => "00010000",
    7185 => "00010000",
    7186 => "00010000",
    7187 => "00010000",
    7188 => "00010000",
    7189 => "00010000",
    7190 => "00010000",
    7191 => "00010000",
    7192 => "00010000",
    7193 => "00010000",
    7194 => "00010000",
    7195 => "00010000",
    7196 => "00010000",
    7197 => "00010000",
    7198 => "00010000",
    7199 => "00010000",
    7200 => "00001111",
    7201 => "00001111",
    7202 => "00001111",
    7203 => "00001111",
    7204 => "00001111",
    7205 => "00001111",
    7206 => "00001111",
    7207 => "00001111",
    7208 => "00001111",
    7209 => "00001111",
    7210 => "00001111",
    7211 => "00001111",
    7212 => "00001111",
    7213 => "00001111",
    7214 => "00001111",
    7215 => "00001111",
    7216 => "00001111",
    7217 => "00001111",
    7218 => "00001111",
    7219 => "00001111",
    7220 => "00001111",
    7221 => "00001111",
    7222 => "00001111",
    7223 => "00001111",
    7224 => "00001111",
    7225 => "00001111",
    7226 => "00001111",
    7227 => "00001111",
    7228 => "00001111",
    7229 => "00001111",
    7230 => "00001111",
    7231 => "00001111",
    7232 => "00001111",
    7233 => "00001111",
    7234 => "00001111",
    7235 => "00001111",
    7236 => "00001111",
    7237 => "00001111",
    7238 => "00001111",
    7239 => "00001111",
    7240 => "00001111",
    7241 => "00001111",
    7242 => "00001111",
    7243 => "00001111",
    7244 => "00001111",
    7245 => "00001111",
    7246 => "00001111",
    7247 => "00001111",
    7248 => "00001111",
    7249 => "00001111",
    7250 => "00001111",
    7251 => "00001111",
    7252 => "00001111",
    7253 => "00001111",
    7254 => "00001111",
    7255 => "00001111",
    7256 => "00001111",
    7257 => "00001111",
    7258 => "00001111",
    7259 => "00001111",
    7260 => "00001111",
    7261 => "00001110",
    7262 => "00001110",
    7263 => "00001110",
    7264 => "00001110",
    7265 => "00001110",
    7266 => "00001110",
    7267 => "00001110",
    7268 => "00001110",
    7269 => "00001110",
    7270 => "00001110",
    7271 => "00001110",
    7272 => "00001110",
    7273 => "00001110",
    7274 => "00001110",
    7275 => "00001110",
    7276 => "00001110",
    7277 => "00001110",
    7278 => "00001110",
    7279 => "00001110",
    7280 => "00001110",
    7281 => "00001110",
    7282 => "00001110",
    7283 => "00001110",
    7284 => "00001110",
    7285 => "00001110",
    7286 => "00001110",
    7287 => "00001110",
    7288 => "00001110",
    7289 => "00001110",
    7290 => "00001110",
    7291 => "00001110",
    7292 => "00001110",
    7293 => "00001110",
    7294 => "00001110",
    7295 => "00001110",
    7296 => "00001110",
    7297 => "00001110",
    7298 => "00001110",
    7299 => "00001110",
    7300 => "00001110",
    7301 => "00001110",
    7302 => "00001110",
    7303 => "00001110",
    7304 => "00001110",
    7305 => "00001110",
    7306 => "00001110",
    7307 => "00001110",
    7308 => "00001110",
    7309 => "00001110",
    7310 => "00001110",
    7311 => "00001110",
    7312 => "00001110",
    7313 => "00001110",
    7314 => "00001110",
    7315 => "00001110",
    7316 => "00001110",
    7317 => "00001110",
    7318 => "00001110",
    7319 => "00001110",
    7320 => "00001110",
    7321 => "00001101",
    7322 => "00001101",
    7323 => "00001101",
    7324 => "00001101",
    7325 => "00001101",
    7326 => "00001101",
    7327 => "00001101",
    7328 => "00001101",
    7329 => "00001101",
    7330 => "00001101",
    7331 => "00001101",
    7332 => "00001101",
    7333 => "00001101",
    7334 => "00001101",
    7335 => "00001101",
    7336 => "00001101",
    7337 => "00001101",
    7338 => "00001101",
    7339 => "00001101",
    7340 => "00001101",
    7341 => "00001101",
    7342 => "00001101",
    7343 => "00001101",
    7344 => "00001101",
    7345 => "00001101",
    7346 => "00001101",
    7347 => "00001101",
    7348 => "00001101",
    7349 => "00001101",
    7350 => "00001101",
    7351 => "00001101",
    7352 => "00001101",
    7353 => "00001101",
    7354 => "00001101",
    7355 => "00001101",
    7356 => "00001101",
    7357 => "00001101",
    7358 => "00001101",
    7359 => "00001101",
    7360 => "00001101",
    7361 => "00001101",
    7362 => "00001101",
    7363 => "00001101",
    7364 => "00001101",
    7365 => "00001101",
    7366 => "00001101",
    7367 => "00001101",
    7368 => "00001101",
    7369 => "00001101",
    7370 => "00001101",
    7371 => "00001101",
    7372 => "00001101",
    7373 => "00001101",
    7374 => "00001101",
    7375 => "00001101",
    7376 => "00001101",
    7377 => "00001101",
    7378 => "00001101",
    7379 => "00001101",
    7380 => "00001101",
    7381 => "00001101",
    7382 => "00001100",
    7383 => "00001100",
    7384 => "00001100",
    7385 => "00001100",
    7386 => "00001100",
    7387 => "00001100",
    7388 => "00001100",
    7389 => "00001100",
    7390 => "00001100",
    7391 => "00001100",
    7392 => "00001100",
    7393 => "00001100",
    7394 => "00001100",
    7395 => "00001100",
    7396 => "00001100",
    7397 => "00001100",
    7398 => "00001100",
    7399 => "00001100",
    7400 => "00001100",
    7401 => "00001100",
    7402 => "00001100",
    7403 => "00001100",
    7404 => "00001100",
    7405 => "00001100",
    7406 => "00001100",
    7407 => "00001100",
    7408 => "00001100",
    7409 => "00001100",
    7410 => "00001100",
    7411 => "00001100",
    7412 => "00001100",
    7413 => "00001100",
    7414 => "00001100",
    7415 => "00001100",
    7416 => "00001100",
    7417 => "00001100",
    7418 => "00001100",
    7419 => "00001100",
    7420 => "00001100",
    7421 => "00001100",
    7422 => "00001100",
    7423 => "00001100",
    7424 => "00001100",
    7425 => "00001100",
    7426 => "00001100",
    7427 => "00001100",
    7428 => "00001100",
    7429 => "00001100",
    7430 => "00001100",
    7431 => "00001100",
    7432 => "00001100",
    7433 => "00001100",
    7434 => "00001100",
    7435 => "00001100",
    7436 => "00001100",
    7437 => "00001100",
    7438 => "00001100",
    7439 => "00001100",
    7440 => "00001100",
    7441 => "00001100",
    7442 => "00001011",
    7443 => "00001011",
    7444 => "00001011",
    7445 => "00001011",
    7446 => "00001011",
    7447 => "00001011",
    7448 => "00001011",
    7449 => "00001011",
    7450 => "00001011",
    7451 => "00001011",
    7452 => "00001011",
    7453 => "00001011",
    7454 => "00001011",
    7455 => "00001011",
    7456 => "00001011",
    7457 => "00001011",
    7458 => "00001011",
    7459 => "00001011",
    7460 => "00001011",
    7461 => "00001011",
    7462 => "00001011",
    7463 => "00001011",
    7464 => "00001011",
    7465 => "00001011",
    7466 => "00001011",
    7467 => "00001011",
    7468 => "00001011",
    7469 => "00001011",
    7470 => "00001011",
    7471 => "00001011",
    7472 => "00001011",
    7473 => "00001011",
    7474 => "00001011",
    7475 => "00001011",
    7476 => "00001011",
    7477 => "00001011",
    7478 => "00001011",
    7479 => "00001011",
    7480 => "00001011",
    7481 => "00001011",
    7482 => "00001011",
    7483 => "00001011",
    7484 => "00001011",
    7485 => "00001011",
    7486 => "00001011",
    7487 => "00001011",
    7488 => "00001011",
    7489 => "00001011",
    7490 => "00001011",
    7491 => "00001011",
    7492 => "00001011",
    7493 => "00001011",
    7494 => "00001011",
    7495 => "00001011",
    7496 => "00001011",
    7497 => "00001011",
    7498 => "00001011",
    7499 => "00001011",
    7500 => "00001011",
    7501 => "00001011",
    7502 => "00001011",
    7503 => "00001011",
    7504 => "00001010",
    7505 => "00001010",
    7506 => "00001010",
    7507 => "00001010",
    7508 => "00001010",
    7509 => "00001010",
    7510 => "00001010",
    7511 => "00001010",
    7512 => "00001010",
    7513 => "00001010",
    7514 => "00001010",
    7515 => "00001010",
    7516 => "00001010",
    7517 => "00001010",
    7518 => "00001010",
    7519 => "00001010",
    7520 => "00001010",
    7521 => "00001010",
    7522 => "00001010",
    7523 => "00001010",
    7524 => "00001010",
    7525 => "00001010",
    7526 => "00001010",
    7527 => "00001010",
    7528 => "00001010",
    7529 => "00001010",
    7530 => "00001010",
    7531 => "00001010",
    7532 => "00001010",
    7533 => "00001010",
    7534 => "00001010",
    7535 => "00001010",
    7536 => "00001010",
    7537 => "00001010",
    7538 => "00001010",
    7539 => "00001010",
    7540 => "00001010",
    7541 => "00001010",
    7542 => "00001010",
    7543 => "00001010",
    7544 => "00001010",
    7545 => "00001010",
    7546 => "00001010",
    7547 => "00001010",
    7548 => "00001010",
    7549 => "00001010",
    7550 => "00001010",
    7551 => "00001010",
    7552 => "00001010",
    7553 => "00001010",
    7554 => "00001010",
    7555 => "00001010",
    7556 => "00001010",
    7557 => "00001010",
    7558 => "00001010",
    7559 => "00001010",
    7560 => "00001010",
    7561 => "00001010",
    7562 => "00001010",
    7563 => "00001010",
    7564 => "00001010",
    7565 => "00001001",
    7566 => "00001001",
    7567 => "00001001",
    7568 => "00001001",
    7569 => "00001001",
    7570 => "00001001",
    7571 => "00001001",
    7572 => "00001001",
    7573 => "00001001",
    7574 => "00001001",
    7575 => "00001001",
    7576 => "00001001",
    7577 => "00001001",
    7578 => "00001001",
    7579 => "00001001",
    7580 => "00001001",
    7581 => "00001001",
    7582 => "00001001",
    7583 => "00001001",
    7584 => "00001001",
    7585 => "00001001",
    7586 => "00001001",
    7587 => "00001001",
    7588 => "00001001",
    7589 => "00001001",
    7590 => "00001001",
    7591 => "00001001",
    7592 => "00001001",
    7593 => "00001001",
    7594 => "00001001",
    7595 => "00001001",
    7596 => "00001001",
    7597 => "00001001",
    7598 => "00001001",
    7599 => "00001001",
    7600 => "00001001",
    7601 => "00001001",
    7602 => "00001001",
    7603 => "00001001",
    7604 => "00001001",
    7605 => "00001001",
    7606 => "00001001",
    7607 => "00001001",
    7608 => "00001001",
    7609 => "00001001",
    7610 => "00001001",
    7611 => "00001001",
    7612 => "00001001",
    7613 => "00001001",
    7614 => "00001001",
    7615 => "00001001",
    7616 => "00001001",
    7617 => "00001001",
    7618 => "00001001",
    7619 => "00001001",
    7620 => "00001001",
    7621 => "00001001",
    7622 => "00001001",
    7623 => "00001001",
    7624 => "00001001",
    7625 => "00001001",
    7626 => "00001001",
    7627 => "00001000",
    7628 => "00001000",
    7629 => "00001000",
    7630 => "00001000",
    7631 => "00001000",
    7632 => "00001000",
    7633 => "00001000",
    7634 => "00001000",
    7635 => "00001000",
    7636 => "00001000",
    7637 => "00001000",
    7638 => "00001000",
    7639 => "00001000",
    7640 => "00001000",
    7641 => "00001000",
    7642 => "00001000",
    7643 => "00001000",
    7644 => "00001000",
    7645 => "00001000",
    7646 => "00001000",
    7647 => "00001000",
    7648 => "00001000",
    7649 => "00001000",
    7650 => "00001000",
    7651 => "00001000",
    7652 => "00001000",
    7653 => "00001000",
    7654 => "00001000",
    7655 => "00001000",
    7656 => "00001000",
    7657 => "00001000",
    7658 => "00001000",
    7659 => "00001000",
    7660 => "00001000",
    7661 => "00001000",
    7662 => "00001000",
    7663 => "00001000",
    7664 => "00001000",
    7665 => "00001000",
    7666 => "00001000",
    7667 => "00001000",
    7668 => "00001000",
    7669 => "00001000",
    7670 => "00001000",
    7671 => "00001000",
    7672 => "00001000",
    7673 => "00001000",
    7674 => "00001000",
    7675 => "00001000",
    7676 => "00001000",
    7677 => "00001000",
    7678 => "00001000",
    7679 => "00001000",
    7680 => "00001000",
    7681 => "00001000",
    7682 => "00001000",
    7683 => "00001000",
    7684 => "00001000",
    7685 => "00001000",
    7686 => "00001000",
    7687 => "00001000",
    7688 => "00000111",
    7689 => "00000111",
    7690 => "00000111",
    7691 => "00000111",
    7692 => "00000111",
    7693 => "00000111",
    7694 => "00000111",
    7695 => "00000111",
    7696 => "00000111",
    7697 => "00000111",
    7698 => "00000111",
    7699 => "00000111",
    7700 => "00000111",
    7701 => "00000111",
    7702 => "00000111",
    7703 => "00000111",
    7704 => "00000111",
    7705 => "00000111",
    7706 => "00000111",
    7707 => "00000111",
    7708 => "00000111",
    7709 => "00000111",
    7710 => "00000111",
    7711 => "00000111",
    7712 => "00000111",
    7713 => "00000111",
    7714 => "00000111",
    7715 => "00000111",
    7716 => "00000111",
    7717 => "00000111",
    7718 => "00000111",
    7719 => "00000111",
    7720 => "00000111",
    7721 => "00000111",
    7722 => "00000111",
    7723 => "00000111",
    7724 => "00000111",
    7725 => "00000111",
    7726 => "00000111",
    7727 => "00000111",
    7728 => "00000111",
    7729 => "00000111",
    7730 => "00000111",
    7731 => "00000111",
    7732 => "00000111",
    7733 => "00000111",
    7734 => "00000111",
    7735 => "00000111",
    7736 => "00000111",
    7737 => "00000111",
    7738 => "00000111",
    7739 => "00000111",
    7740 => "00000111",
    7741 => "00000111",
    7742 => "00000111",
    7743 => "00000111",
    7744 => "00000111",
    7745 => "00000111",
    7746 => "00000111",
    7747 => "00000111",
    7748 => "00000111",
    7749 => "00000111",
    7750 => "00000111",
    7751 => "00000110",
    7752 => "00000110",
    7753 => "00000110",
    7754 => "00000110",
    7755 => "00000110",
    7756 => "00000110",
    7757 => "00000110",
    7758 => "00000110",
    7759 => "00000110",
    7760 => "00000110",
    7761 => "00000110",
    7762 => "00000110",
    7763 => "00000110",
    7764 => "00000110",
    7765 => "00000110",
    7766 => "00000110",
    7767 => "00000110",
    7768 => "00000110",
    7769 => "00000110",
    7770 => "00000110",
    7771 => "00000110",
    7772 => "00000110",
    7773 => "00000110",
    7774 => "00000110",
    7775 => "00000110",
    7776 => "00000110",
    7777 => "00000110",
    7778 => "00000110",
    7779 => "00000110",
    7780 => "00000110",
    7781 => "00000110",
    7782 => "00000110",
    7783 => "00000110",
    7784 => "00000110",
    7785 => "00000110",
    7786 => "00000110",
    7787 => "00000110",
    7788 => "00000110",
    7789 => "00000110",
    7790 => "00000110",
    7791 => "00000110",
    7792 => "00000110",
    7793 => "00000110",
    7794 => "00000110",
    7795 => "00000110",
    7796 => "00000110",
    7797 => "00000110",
    7798 => "00000110",
    7799 => "00000110",
    7800 => "00000110",
    7801 => "00000110",
    7802 => "00000110",
    7803 => "00000110",
    7804 => "00000110",
    7805 => "00000110",
    7806 => "00000110",
    7807 => "00000110",
    7808 => "00000110",
    7809 => "00000110",
    7810 => "00000110",
    7811 => "00000110",
    7812 => "00000110",
    7813 => "00000101",
    7814 => "00000101",
    7815 => "00000101",
    7816 => "00000101",
    7817 => "00000101",
    7818 => "00000101",
    7819 => "00000101",
    7820 => "00000101",
    7821 => "00000101",
    7822 => "00000101",
    7823 => "00000101",
    7824 => "00000101",
    7825 => "00000101",
    7826 => "00000101",
    7827 => "00000101",
    7828 => "00000101",
    7829 => "00000101",
    7830 => "00000101",
    7831 => "00000101",
    7832 => "00000101",
    7833 => "00000101",
    7834 => "00000101",
    7835 => "00000101",
    7836 => "00000101",
    7837 => "00000101",
    7838 => "00000101",
    7839 => "00000101",
    7840 => "00000101",
    7841 => "00000101",
    7842 => "00000101",
    7843 => "00000101",
    7844 => "00000101",
    7845 => "00000101",
    7846 => "00000101",
    7847 => "00000101",
    7848 => "00000101",
    7849 => "00000101",
    7850 => "00000101",
    7851 => "00000101",
    7852 => "00000101",
    7853 => "00000101",
    7854 => "00000101",
    7855 => "00000101",
    7856 => "00000101",
    7857 => "00000101",
    7858 => "00000101",
    7859 => "00000101",
    7860 => "00000101",
    7861 => "00000101",
    7862 => "00000101",
    7863 => "00000101",
    7864 => "00000101",
    7865 => "00000101",
    7866 => "00000101",
    7867 => "00000101",
    7868 => "00000101",
    7869 => "00000101",
    7870 => "00000101",
    7871 => "00000101",
    7872 => "00000101",
    7873 => "00000101",
    7874 => "00000101",
    7875 => "00000101",
    7876 => "00000100",
    7877 => "00000100",
    7878 => "00000100",
    7879 => "00000100",
    7880 => "00000100",
    7881 => "00000100",
    7882 => "00000100",
    7883 => "00000100",
    7884 => "00000100",
    7885 => "00000100",
    7886 => "00000100",
    7887 => "00000100",
    7888 => "00000100",
    7889 => "00000100",
    7890 => "00000100",
    7891 => "00000100",
    7892 => "00000100",
    7893 => "00000100",
    7894 => "00000100",
    7895 => "00000100",
    7896 => "00000100",
    7897 => "00000100",
    7898 => "00000100",
    7899 => "00000100",
    7900 => "00000100",
    7901 => "00000100",
    7902 => "00000100",
    7903 => "00000100",
    7904 => "00000100",
    7905 => "00000100",
    7906 => "00000100",
    7907 => "00000100",
    7908 => "00000100",
    7909 => "00000100",
    7910 => "00000100",
    7911 => "00000100",
    7912 => "00000100",
    7913 => "00000100",
    7914 => "00000100",
    7915 => "00000100",
    7916 => "00000100",
    7917 => "00000100",
    7918 => "00000100",
    7919 => "00000100",
    7920 => "00000100",
    7921 => "00000100",
    7922 => "00000100",
    7923 => "00000100",
    7924 => "00000100",
    7925 => "00000100",
    7926 => "00000100",
    7927 => "00000100",
    7928 => "00000100",
    7929 => "00000100",
    7930 => "00000100",
    7931 => "00000100",
    7932 => "00000100",
    7933 => "00000100",
    7934 => "00000100",
    7935 => "00000100",
    7936 => "00000100",
    7937 => "00000100",
    7938 => "00000011",
    7939 => "00000011",
    7940 => "00000011",
    7941 => "00000011",
    7942 => "00000011",
    7943 => "00000011",
    7944 => "00000011",
    7945 => "00000011",
    7946 => "00000011",
    7947 => "00000011",
    7948 => "00000011",
    7949 => "00000011",
    7950 => "00000011",
    7951 => "00000011",
    7952 => "00000011",
    7953 => "00000011",
    7954 => "00000011",
    7955 => "00000011",
    7956 => "00000011",
    7957 => "00000011",
    7958 => "00000011",
    7959 => "00000011",
    7960 => "00000011",
    7961 => "00000011",
    7962 => "00000011",
    7963 => "00000011",
    7964 => "00000011",
    7965 => "00000011",
    7966 => "00000011",
    7967 => "00000011",
    7968 => "00000011",
    7969 => "00000011",
    7970 => "00000011",
    7971 => "00000011",
    7972 => "00000011",
    7973 => "00000011",
    7974 => "00000011",
    7975 => "00000011",
    7976 => "00000011",
    7977 => "00000011",
    7978 => "00000011",
    7979 => "00000011",
    7980 => "00000011",
    7981 => "00000011",
    7982 => "00000011",
    7983 => "00000011",
    7984 => "00000011",
    7985 => "00000011",
    7986 => "00000011",
    7987 => "00000011",
    7988 => "00000011",
    7989 => "00000011",
    7990 => "00000011",
    7991 => "00000011",
    7992 => "00000011",
    7993 => "00000011",
    7994 => "00000011",
    7995 => "00000011",
    7996 => "00000011",
    7997 => "00000011",
    7998 => "00000011",
    7999 => "00000011",
    8000 => "00000011",
    8001 => "00000011",
    8002 => "00000010",
    8003 => "00000010",
    8004 => "00000010",
    8005 => "00000010",
    8006 => "00000010",
    8007 => "00000010",
    8008 => "00000010",
    8009 => "00000010",
    8010 => "00000010",
    8011 => "00000010",
    8012 => "00000010",
    8013 => "00000010",
    8014 => "00000010",
    8015 => "00000010",
    8016 => "00000010",
    8017 => "00000010",
    8018 => "00000010",
    8019 => "00000010",
    8020 => "00000010",
    8021 => "00000010",
    8022 => "00000010",
    8023 => "00000010",
    8024 => "00000010",
    8025 => "00000010",
    8026 => "00000010",
    8027 => "00000010",
    8028 => "00000010",
    8029 => "00000010",
    8030 => "00000010",
    8031 => "00000010",
    8032 => "00000010",
    8033 => "00000010",
    8034 => "00000010",
    8035 => "00000010",
    8036 => "00000010",
    8037 => "00000010",
    8038 => "00000010",
    8039 => "00000010",
    8040 => "00000010",
    8041 => "00000010",
    8042 => "00000010",
    8043 => "00000010",
    8044 => "00000010",
    8045 => "00000010",
    8046 => "00000010",
    8047 => "00000010",
    8048 => "00000010",
    8049 => "00000010",
    8050 => "00000010",
    8051 => "00000010",
    8052 => "00000010",
    8053 => "00000010",
    8054 => "00000010",
    8055 => "00000010",
    8056 => "00000010",
    8057 => "00000010",
    8058 => "00000010",
    8059 => "00000010",
    8060 => "00000010",
    8061 => "00000010",
    8062 => "00000010",
    8063 => "00000010",
    8064 => "00000010",
    8065 => "00000001",
    8066 => "00000001",
    8067 => "00000001",
    8068 => "00000001",
    8069 => "00000001",
    8070 => "00000001",
    8071 => "00000001",
    8072 => "00000001",
    8073 => "00000001",
    8074 => "00000001",
    8075 => "00000001",
    8076 => "00000001",
    8077 => "00000001",
    8078 => "00000001",
    8079 => "00000001",
    8080 => "00000001",
    8081 => "00000001",
    8082 => "00000001",
    8083 => "00000001",
    8084 => "00000001",
    8085 => "00000001",
    8086 => "00000001",
    8087 => "00000001",
    8088 => "00000001",
    8089 => "00000001",
    8090 => "00000001",
    8091 => "00000001",
    8092 => "00000001",
    8093 => "00000001",
    8094 => "00000001",
    8095 => "00000001",
    8096 => "00000001",
    8097 => "00000001",
    8098 => "00000001",
    8099 => "00000001",
    8100 => "00000001",
    8101 => "00000001",
    8102 => "00000001",
    8103 => "00000001",
    8104 => "00000001",
    8105 => "00000001",
    8106 => "00000001",
    8107 => "00000001",
    8108 => "00000001",
    8109 => "00000001",
    8110 => "00000001",
    8111 => "00000001",
    8112 => "00000001",
    8113 => "00000001",
    8114 => "00000001",
    8115 => "00000001",
    8116 => "00000001",
    8117 => "00000001",
    8118 => "00000001",
    8119 => "00000001",
    8120 => "00000001",
    8121 => "00000001",
    8122 => "00000001",
    8123 => "00000001",
    8124 => "00000001",
    8125 => "00000001",
    8126 => "00000001",
    8127 => "00000001",
    8128 => "00000001",
    8129 => "00000000",
    8130 => "00000000",
    8131 => "00000000",
    8132 => "00000000",
    8133 => "00000000",
    8134 => "00000000",
    8135 => "00000000",
    8136 => "00000000",
    8137 => "00000000",
    8138 => "00000000",
    8139 => "00000000",
    8140 => "00000000",
    8141 => "00000000",
    8142 => "00000000",
    8143 => "00000000",
    8144 => "00000000",
    8145 => "00000000",
    8146 => "00000000",
    8147 => "00000000",
    8148 => "00000000",
    8149 => "00000000",
    8150 => "00000000",
    8151 => "00000000",
    8152 => "00000000",
    8153 => "00000000",
    8154 => "00000000",
    8155 => "00000000",
    8156 => "00000000",
    8157 => "00000000",
    8158 => "00000000",
    8159 => "00000000",
    8160 => "00000000",
    8161 => "00000000",
    8162 => "00000000",
    8163 => "00000000",
    8164 => "00000000",
    8165 => "00000000",
    8166 => "00000000",
    8167 => "00000000",
    8168 => "00000000",
    8169 => "00000000",
    8170 => "00000000",
    8171 => "00000000",
    8172 => "00000000",
    8173 => "00000000",
    8174 => "00000000",
    8175 => "00000000",
    8176 => "00000000",
    8177 => "00000000",
    8178 => "00000000",
    8179 => "00000000",
    8180 => "00000000",
    8181 => "00000000",
    8182 => "00000000",
    8183 => "00000000",
    8184 => "00000000",
    8185 => "00000000",
    8186 => "00000000",
    8187 => "00000000",
    8188 => "00000000",
    8189 => "00000000",
    8190 => "00000000",
    8191 => "00000000");
  signal q_unbuf : std_logic_vector(7 downto 0);
begin
   process (address)
   begin
     case address is
      when "0000000000000" => q_unbuf <= my_rom(0);
      when "0000000000001" => q_unbuf <= my_rom(1);
      when "0000000000010" => q_unbuf <= my_rom(2);
      when "0000000000011" => q_unbuf <= my_rom(3);
      when "0000000000100" => q_unbuf <= my_rom(4);
      when "0000000000101" => q_unbuf <= my_rom(5);
      when "0000000000110" => q_unbuf <= my_rom(6);
      when "0000000000111" => q_unbuf <= my_rom(7);
      when "0000000001000" => q_unbuf <= my_rom(8);
      when "0000000001001" => q_unbuf <= my_rom(9);
      when "0000000001010" => q_unbuf <= my_rom(10);
      when "0000000001011" => q_unbuf <= my_rom(11);
      when "0000000001100" => q_unbuf <= my_rom(12);
      when "0000000001101" => q_unbuf <= my_rom(13);
      when "0000000001110" => q_unbuf <= my_rom(14);
      when "0000000001111" => q_unbuf <= my_rom(15);
      when "0000000010000" => q_unbuf <= my_rom(16);
      when "0000000010001" => q_unbuf <= my_rom(17);
      when "0000000010010" => q_unbuf <= my_rom(18);
      when "0000000010011" => q_unbuf <= my_rom(19);
      when "0000000010100" => q_unbuf <= my_rom(20);
      when "0000000010101" => q_unbuf <= my_rom(21);
      when "0000000010110" => q_unbuf <= my_rom(22);
      when "0000000010111" => q_unbuf <= my_rom(23);
      when "0000000011000" => q_unbuf <= my_rom(24);
      when "0000000011001" => q_unbuf <= my_rom(25);
      when "0000000011010" => q_unbuf <= my_rom(26);
      when "0000000011011" => q_unbuf <= my_rom(27);
      when "0000000011100" => q_unbuf <= my_rom(28);
      when "0000000011101" => q_unbuf <= my_rom(29);
      when "0000000011110" => q_unbuf <= my_rom(30);
      when "0000000011111" => q_unbuf <= my_rom(31);
      when "0000000100000" => q_unbuf <= my_rom(32);
      when "0000000100001" => q_unbuf <= my_rom(33);
      when "0000000100010" => q_unbuf <= my_rom(34);
      when "0000000100011" => q_unbuf <= my_rom(35);
      when "0000000100100" => q_unbuf <= my_rom(36);
      when "0000000100101" => q_unbuf <= my_rom(37);
      when "0000000100110" => q_unbuf <= my_rom(38);
      when "0000000100111" => q_unbuf <= my_rom(39);
      when "0000000101000" => q_unbuf <= my_rom(40);
      when "0000000101001" => q_unbuf <= my_rom(41);
      when "0000000101010" => q_unbuf <= my_rom(42);
      when "0000000101011" => q_unbuf <= my_rom(43);
      when "0000000101100" => q_unbuf <= my_rom(44);
      when "0000000101101" => q_unbuf <= my_rom(45);
      when "0000000101110" => q_unbuf <= my_rom(46);
      when "0000000101111" => q_unbuf <= my_rom(47);
      when "0000000110000" => q_unbuf <= my_rom(48);
      when "0000000110001" => q_unbuf <= my_rom(49);
      when "0000000110010" => q_unbuf <= my_rom(50);
      when "0000000110011" => q_unbuf <= my_rom(51);
      when "0000000110100" => q_unbuf <= my_rom(52);
      when "0000000110101" => q_unbuf <= my_rom(53);
      when "0000000110110" => q_unbuf <= my_rom(54);
      when "0000000110111" => q_unbuf <= my_rom(55);
      when "0000000111000" => q_unbuf <= my_rom(56);
      when "0000000111001" => q_unbuf <= my_rom(57);
      when "0000000111010" => q_unbuf <= my_rom(58);
      when "0000000111011" => q_unbuf <= my_rom(59);
      when "0000000111100" => q_unbuf <= my_rom(60);
      when "0000000111101" => q_unbuf <= my_rom(61);
      when "0000000111110" => q_unbuf <= my_rom(62);
      when "0000000111111" => q_unbuf <= my_rom(63);
      when "0000001000000" => q_unbuf <= my_rom(64);
      when "0000001000001" => q_unbuf <= my_rom(65);
      when "0000001000010" => q_unbuf <= my_rom(66);
      when "0000001000011" => q_unbuf <= my_rom(67);
      when "0000001000100" => q_unbuf <= my_rom(68);
      when "0000001000101" => q_unbuf <= my_rom(69);
      when "0000001000110" => q_unbuf <= my_rom(70);
      when "0000001000111" => q_unbuf <= my_rom(71);
      when "0000001001000" => q_unbuf <= my_rom(72);
      when "0000001001001" => q_unbuf <= my_rom(73);
      when "0000001001010" => q_unbuf <= my_rom(74);
      when "0000001001011" => q_unbuf <= my_rom(75);
      when "0000001001100" => q_unbuf <= my_rom(76);
      when "0000001001101" => q_unbuf <= my_rom(77);
      when "0000001001110" => q_unbuf <= my_rom(78);
      when "0000001001111" => q_unbuf <= my_rom(79);
      when "0000001010000" => q_unbuf <= my_rom(80);
      when "0000001010001" => q_unbuf <= my_rom(81);
      when "0000001010010" => q_unbuf <= my_rom(82);
      when "0000001010011" => q_unbuf <= my_rom(83);
      when "0000001010100" => q_unbuf <= my_rom(84);
      when "0000001010101" => q_unbuf <= my_rom(85);
      when "0000001010110" => q_unbuf <= my_rom(86);
      when "0000001010111" => q_unbuf <= my_rom(87);
      when "0000001011000" => q_unbuf <= my_rom(88);
      when "0000001011001" => q_unbuf <= my_rom(89);
      when "0000001011010" => q_unbuf <= my_rom(90);
      when "0000001011011" => q_unbuf <= my_rom(91);
      when "0000001011100" => q_unbuf <= my_rom(92);
      when "0000001011101" => q_unbuf <= my_rom(93);
      when "0000001011110" => q_unbuf <= my_rom(94);
      when "0000001011111" => q_unbuf <= my_rom(95);
      when "0000001100000" => q_unbuf <= my_rom(96);
      when "0000001100001" => q_unbuf <= my_rom(97);
      when "0000001100010" => q_unbuf <= my_rom(98);
      when "0000001100011" => q_unbuf <= my_rom(99);
      when "0000001100100" => q_unbuf <= my_rom(100);
      when "0000001100101" => q_unbuf <= my_rom(101);
      when "0000001100110" => q_unbuf <= my_rom(102);
      when "0000001100111" => q_unbuf <= my_rom(103);
      when "0000001101000" => q_unbuf <= my_rom(104);
      when "0000001101001" => q_unbuf <= my_rom(105);
      when "0000001101010" => q_unbuf <= my_rom(106);
      when "0000001101011" => q_unbuf <= my_rom(107);
      when "0000001101100" => q_unbuf <= my_rom(108);
      when "0000001101101" => q_unbuf <= my_rom(109);
      when "0000001101110" => q_unbuf <= my_rom(110);
      when "0000001101111" => q_unbuf <= my_rom(111);
      when "0000001110000" => q_unbuf <= my_rom(112);
      when "0000001110001" => q_unbuf <= my_rom(113);
      when "0000001110010" => q_unbuf <= my_rom(114);
      when "0000001110011" => q_unbuf <= my_rom(115);
      when "0000001110100" => q_unbuf <= my_rom(116);
      when "0000001110101" => q_unbuf <= my_rom(117);
      when "0000001110110" => q_unbuf <= my_rom(118);
      when "0000001110111" => q_unbuf <= my_rom(119);
      when "0000001111000" => q_unbuf <= my_rom(120);
      when "0000001111001" => q_unbuf <= my_rom(121);
      when "0000001111010" => q_unbuf <= my_rom(122);
      when "0000001111011" => q_unbuf <= my_rom(123);
      when "0000001111100" => q_unbuf <= my_rom(124);
      when "0000001111101" => q_unbuf <= my_rom(125);
      when "0000001111110" => q_unbuf <= my_rom(126);
      when "0000001111111" => q_unbuf <= my_rom(127);
      when "0000010000000" => q_unbuf <= my_rom(128);
      when "0000010000001" => q_unbuf <= my_rom(129);
      when "0000010000010" => q_unbuf <= my_rom(130);
      when "0000010000011" => q_unbuf <= my_rom(131);
      when "0000010000100" => q_unbuf <= my_rom(132);
      when "0000010000101" => q_unbuf <= my_rom(133);
      when "0000010000110" => q_unbuf <= my_rom(134);
      when "0000010000111" => q_unbuf <= my_rom(135);
      when "0000010001000" => q_unbuf <= my_rom(136);
      when "0000010001001" => q_unbuf <= my_rom(137);
      when "0000010001010" => q_unbuf <= my_rom(138);
      when "0000010001011" => q_unbuf <= my_rom(139);
      when "0000010001100" => q_unbuf <= my_rom(140);
      when "0000010001101" => q_unbuf <= my_rom(141);
      when "0000010001110" => q_unbuf <= my_rom(142);
      when "0000010001111" => q_unbuf <= my_rom(143);
      when "0000010010000" => q_unbuf <= my_rom(144);
      when "0000010010001" => q_unbuf <= my_rom(145);
      when "0000010010010" => q_unbuf <= my_rom(146);
      when "0000010010011" => q_unbuf <= my_rom(147);
      when "0000010010100" => q_unbuf <= my_rom(148);
      when "0000010010101" => q_unbuf <= my_rom(149);
      when "0000010010110" => q_unbuf <= my_rom(150);
      when "0000010010111" => q_unbuf <= my_rom(151);
      when "0000010011000" => q_unbuf <= my_rom(152);
      when "0000010011001" => q_unbuf <= my_rom(153);
      when "0000010011010" => q_unbuf <= my_rom(154);
      when "0000010011011" => q_unbuf <= my_rom(155);
      when "0000010011100" => q_unbuf <= my_rom(156);
      when "0000010011101" => q_unbuf <= my_rom(157);
      when "0000010011110" => q_unbuf <= my_rom(158);
      when "0000010011111" => q_unbuf <= my_rom(159);
      when "0000010100000" => q_unbuf <= my_rom(160);
      when "0000010100001" => q_unbuf <= my_rom(161);
      when "0000010100010" => q_unbuf <= my_rom(162);
      when "0000010100011" => q_unbuf <= my_rom(163);
      when "0000010100100" => q_unbuf <= my_rom(164);
      when "0000010100101" => q_unbuf <= my_rom(165);
      when "0000010100110" => q_unbuf <= my_rom(166);
      when "0000010100111" => q_unbuf <= my_rom(167);
      when "0000010101000" => q_unbuf <= my_rom(168);
      when "0000010101001" => q_unbuf <= my_rom(169);
      when "0000010101010" => q_unbuf <= my_rom(170);
      when "0000010101011" => q_unbuf <= my_rom(171);
      when "0000010101100" => q_unbuf <= my_rom(172);
      when "0000010101101" => q_unbuf <= my_rom(173);
      when "0000010101110" => q_unbuf <= my_rom(174);
      when "0000010101111" => q_unbuf <= my_rom(175);
      when "0000010110000" => q_unbuf <= my_rom(176);
      when "0000010110001" => q_unbuf <= my_rom(177);
      when "0000010110010" => q_unbuf <= my_rom(178);
      when "0000010110011" => q_unbuf <= my_rom(179);
      when "0000010110100" => q_unbuf <= my_rom(180);
      when "0000010110101" => q_unbuf <= my_rom(181);
      when "0000010110110" => q_unbuf <= my_rom(182);
      when "0000010110111" => q_unbuf <= my_rom(183);
      when "0000010111000" => q_unbuf <= my_rom(184);
      when "0000010111001" => q_unbuf <= my_rom(185);
      when "0000010111010" => q_unbuf <= my_rom(186);
      when "0000010111011" => q_unbuf <= my_rom(187);
      when "0000010111100" => q_unbuf <= my_rom(188);
      when "0000010111101" => q_unbuf <= my_rom(189);
      when "0000010111110" => q_unbuf <= my_rom(190);
      when "0000010111111" => q_unbuf <= my_rom(191);
      when "0000011000000" => q_unbuf <= my_rom(192);
      when "0000011000001" => q_unbuf <= my_rom(193);
      when "0000011000010" => q_unbuf <= my_rom(194);
      when "0000011000011" => q_unbuf <= my_rom(195);
      when "0000011000100" => q_unbuf <= my_rom(196);
      when "0000011000101" => q_unbuf <= my_rom(197);
      when "0000011000110" => q_unbuf <= my_rom(198);
      when "0000011000111" => q_unbuf <= my_rom(199);
      when "0000011001000" => q_unbuf <= my_rom(200);
      when "0000011001001" => q_unbuf <= my_rom(201);
      when "0000011001010" => q_unbuf <= my_rom(202);
      when "0000011001011" => q_unbuf <= my_rom(203);
      when "0000011001100" => q_unbuf <= my_rom(204);
      when "0000011001101" => q_unbuf <= my_rom(205);
      when "0000011001110" => q_unbuf <= my_rom(206);
      when "0000011001111" => q_unbuf <= my_rom(207);
      when "0000011010000" => q_unbuf <= my_rom(208);
      when "0000011010001" => q_unbuf <= my_rom(209);
      when "0000011010010" => q_unbuf <= my_rom(210);
      when "0000011010011" => q_unbuf <= my_rom(211);
      when "0000011010100" => q_unbuf <= my_rom(212);
      when "0000011010101" => q_unbuf <= my_rom(213);
      when "0000011010110" => q_unbuf <= my_rom(214);
      when "0000011010111" => q_unbuf <= my_rom(215);
      when "0000011011000" => q_unbuf <= my_rom(216);
      when "0000011011001" => q_unbuf <= my_rom(217);
      when "0000011011010" => q_unbuf <= my_rom(218);
      when "0000011011011" => q_unbuf <= my_rom(219);
      when "0000011011100" => q_unbuf <= my_rom(220);
      when "0000011011101" => q_unbuf <= my_rom(221);
      when "0000011011110" => q_unbuf <= my_rom(222);
      when "0000011011111" => q_unbuf <= my_rom(223);
      when "0000011100000" => q_unbuf <= my_rom(224);
      when "0000011100001" => q_unbuf <= my_rom(225);
      when "0000011100010" => q_unbuf <= my_rom(226);
      when "0000011100011" => q_unbuf <= my_rom(227);
      when "0000011100100" => q_unbuf <= my_rom(228);
      when "0000011100101" => q_unbuf <= my_rom(229);
      when "0000011100110" => q_unbuf <= my_rom(230);
      when "0000011100111" => q_unbuf <= my_rom(231);
      when "0000011101000" => q_unbuf <= my_rom(232);
      when "0000011101001" => q_unbuf <= my_rom(233);
      when "0000011101010" => q_unbuf <= my_rom(234);
      when "0000011101011" => q_unbuf <= my_rom(235);
      when "0000011101100" => q_unbuf <= my_rom(236);
      when "0000011101101" => q_unbuf <= my_rom(237);
      when "0000011101110" => q_unbuf <= my_rom(238);
      when "0000011101111" => q_unbuf <= my_rom(239);
      when "0000011110000" => q_unbuf <= my_rom(240);
      when "0000011110001" => q_unbuf <= my_rom(241);
      when "0000011110010" => q_unbuf <= my_rom(242);
      when "0000011110011" => q_unbuf <= my_rom(243);
      when "0000011110100" => q_unbuf <= my_rom(244);
      when "0000011110101" => q_unbuf <= my_rom(245);
      when "0000011110110" => q_unbuf <= my_rom(246);
      when "0000011110111" => q_unbuf <= my_rom(247);
      when "0000011111000" => q_unbuf <= my_rom(248);
      when "0000011111001" => q_unbuf <= my_rom(249);
      when "0000011111010" => q_unbuf <= my_rom(250);
      when "0000011111011" => q_unbuf <= my_rom(251);
      when "0000011111100" => q_unbuf <= my_rom(252);
      when "0000011111101" => q_unbuf <= my_rom(253);
      when "0000011111110" => q_unbuf <= my_rom(254);
      when "0000011111111" => q_unbuf <= my_rom(255);
      when "0000100000000" => q_unbuf <= my_rom(256);
      when "0000100000001" => q_unbuf <= my_rom(257);
      when "0000100000010" => q_unbuf <= my_rom(258);
      when "0000100000011" => q_unbuf <= my_rom(259);
      when "0000100000100" => q_unbuf <= my_rom(260);
      when "0000100000101" => q_unbuf <= my_rom(261);
      when "0000100000110" => q_unbuf <= my_rom(262);
      when "0000100000111" => q_unbuf <= my_rom(263);
      when "0000100001000" => q_unbuf <= my_rom(264);
      when "0000100001001" => q_unbuf <= my_rom(265);
      when "0000100001010" => q_unbuf <= my_rom(266);
      when "0000100001011" => q_unbuf <= my_rom(267);
      when "0000100001100" => q_unbuf <= my_rom(268);
      when "0000100001101" => q_unbuf <= my_rom(269);
      when "0000100001110" => q_unbuf <= my_rom(270);
      when "0000100001111" => q_unbuf <= my_rom(271);
      when "0000100010000" => q_unbuf <= my_rom(272);
      when "0000100010001" => q_unbuf <= my_rom(273);
      when "0000100010010" => q_unbuf <= my_rom(274);
      when "0000100010011" => q_unbuf <= my_rom(275);
      when "0000100010100" => q_unbuf <= my_rom(276);
      when "0000100010101" => q_unbuf <= my_rom(277);
      when "0000100010110" => q_unbuf <= my_rom(278);
      when "0000100010111" => q_unbuf <= my_rom(279);
      when "0000100011000" => q_unbuf <= my_rom(280);
      when "0000100011001" => q_unbuf <= my_rom(281);
      when "0000100011010" => q_unbuf <= my_rom(282);
      when "0000100011011" => q_unbuf <= my_rom(283);
      when "0000100011100" => q_unbuf <= my_rom(284);
      when "0000100011101" => q_unbuf <= my_rom(285);
      when "0000100011110" => q_unbuf <= my_rom(286);
      when "0000100011111" => q_unbuf <= my_rom(287);
      when "0000100100000" => q_unbuf <= my_rom(288);
      when "0000100100001" => q_unbuf <= my_rom(289);
      when "0000100100010" => q_unbuf <= my_rom(290);
      when "0000100100011" => q_unbuf <= my_rom(291);
      when "0000100100100" => q_unbuf <= my_rom(292);
      when "0000100100101" => q_unbuf <= my_rom(293);
      when "0000100100110" => q_unbuf <= my_rom(294);
      when "0000100100111" => q_unbuf <= my_rom(295);
      when "0000100101000" => q_unbuf <= my_rom(296);
      when "0000100101001" => q_unbuf <= my_rom(297);
      when "0000100101010" => q_unbuf <= my_rom(298);
      when "0000100101011" => q_unbuf <= my_rom(299);
      when "0000100101100" => q_unbuf <= my_rom(300);
      when "0000100101101" => q_unbuf <= my_rom(301);
      when "0000100101110" => q_unbuf <= my_rom(302);
      when "0000100101111" => q_unbuf <= my_rom(303);
      when "0000100110000" => q_unbuf <= my_rom(304);
      when "0000100110001" => q_unbuf <= my_rom(305);
      when "0000100110010" => q_unbuf <= my_rom(306);
      when "0000100110011" => q_unbuf <= my_rom(307);
      when "0000100110100" => q_unbuf <= my_rom(308);
      when "0000100110101" => q_unbuf <= my_rom(309);
      when "0000100110110" => q_unbuf <= my_rom(310);
      when "0000100110111" => q_unbuf <= my_rom(311);
      when "0000100111000" => q_unbuf <= my_rom(312);
      when "0000100111001" => q_unbuf <= my_rom(313);
      when "0000100111010" => q_unbuf <= my_rom(314);
      when "0000100111011" => q_unbuf <= my_rom(315);
      when "0000100111100" => q_unbuf <= my_rom(316);
      when "0000100111101" => q_unbuf <= my_rom(317);
      when "0000100111110" => q_unbuf <= my_rom(318);
      when "0000100111111" => q_unbuf <= my_rom(319);
      when "0000101000000" => q_unbuf <= my_rom(320);
      when "0000101000001" => q_unbuf <= my_rom(321);
      when "0000101000010" => q_unbuf <= my_rom(322);
      when "0000101000011" => q_unbuf <= my_rom(323);
      when "0000101000100" => q_unbuf <= my_rom(324);
      when "0000101000101" => q_unbuf <= my_rom(325);
      when "0000101000110" => q_unbuf <= my_rom(326);
      when "0000101000111" => q_unbuf <= my_rom(327);
      when "0000101001000" => q_unbuf <= my_rom(328);
      when "0000101001001" => q_unbuf <= my_rom(329);
      when "0000101001010" => q_unbuf <= my_rom(330);
      when "0000101001011" => q_unbuf <= my_rom(331);
      when "0000101001100" => q_unbuf <= my_rom(332);
      when "0000101001101" => q_unbuf <= my_rom(333);
      when "0000101001110" => q_unbuf <= my_rom(334);
      when "0000101001111" => q_unbuf <= my_rom(335);
      when "0000101010000" => q_unbuf <= my_rom(336);
      when "0000101010001" => q_unbuf <= my_rom(337);
      when "0000101010010" => q_unbuf <= my_rom(338);
      when "0000101010011" => q_unbuf <= my_rom(339);
      when "0000101010100" => q_unbuf <= my_rom(340);
      when "0000101010101" => q_unbuf <= my_rom(341);
      when "0000101010110" => q_unbuf <= my_rom(342);
      when "0000101010111" => q_unbuf <= my_rom(343);
      when "0000101011000" => q_unbuf <= my_rom(344);
      when "0000101011001" => q_unbuf <= my_rom(345);
      when "0000101011010" => q_unbuf <= my_rom(346);
      when "0000101011011" => q_unbuf <= my_rom(347);
      when "0000101011100" => q_unbuf <= my_rom(348);
      when "0000101011101" => q_unbuf <= my_rom(349);
      when "0000101011110" => q_unbuf <= my_rom(350);
      when "0000101011111" => q_unbuf <= my_rom(351);
      when "0000101100000" => q_unbuf <= my_rom(352);
      when "0000101100001" => q_unbuf <= my_rom(353);
      when "0000101100010" => q_unbuf <= my_rom(354);
      when "0000101100011" => q_unbuf <= my_rom(355);
      when "0000101100100" => q_unbuf <= my_rom(356);
      when "0000101100101" => q_unbuf <= my_rom(357);
      when "0000101100110" => q_unbuf <= my_rom(358);
      when "0000101100111" => q_unbuf <= my_rom(359);
      when "0000101101000" => q_unbuf <= my_rom(360);
      when "0000101101001" => q_unbuf <= my_rom(361);
      when "0000101101010" => q_unbuf <= my_rom(362);
      when "0000101101011" => q_unbuf <= my_rom(363);
      when "0000101101100" => q_unbuf <= my_rom(364);
      when "0000101101101" => q_unbuf <= my_rom(365);
      when "0000101101110" => q_unbuf <= my_rom(366);
      when "0000101101111" => q_unbuf <= my_rom(367);
      when "0000101110000" => q_unbuf <= my_rom(368);
      when "0000101110001" => q_unbuf <= my_rom(369);
      when "0000101110010" => q_unbuf <= my_rom(370);
      when "0000101110011" => q_unbuf <= my_rom(371);
      when "0000101110100" => q_unbuf <= my_rom(372);
      when "0000101110101" => q_unbuf <= my_rom(373);
      when "0000101110110" => q_unbuf <= my_rom(374);
      when "0000101110111" => q_unbuf <= my_rom(375);
      when "0000101111000" => q_unbuf <= my_rom(376);
      when "0000101111001" => q_unbuf <= my_rom(377);
      when "0000101111010" => q_unbuf <= my_rom(378);
      when "0000101111011" => q_unbuf <= my_rom(379);
      when "0000101111100" => q_unbuf <= my_rom(380);
      when "0000101111101" => q_unbuf <= my_rom(381);
      when "0000101111110" => q_unbuf <= my_rom(382);
      when "0000101111111" => q_unbuf <= my_rom(383);
      when "0000110000000" => q_unbuf <= my_rom(384);
      when "0000110000001" => q_unbuf <= my_rom(385);
      when "0000110000010" => q_unbuf <= my_rom(386);
      when "0000110000011" => q_unbuf <= my_rom(387);
      when "0000110000100" => q_unbuf <= my_rom(388);
      when "0000110000101" => q_unbuf <= my_rom(389);
      when "0000110000110" => q_unbuf <= my_rom(390);
      when "0000110000111" => q_unbuf <= my_rom(391);
      when "0000110001000" => q_unbuf <= my_rom(392);
      when "0000110001001" => q_unbuf <= my_rom(393);
      when "0000110001010" => q_unbuf <= my_rom(394);
      when "0000110001011" => q_unbuf <= my_rom(395);
      when "0000110001100" => q_unbuf <= my_rom(396);
      when "0000110001101" => q_unbuf <= my_rom(397);
      when "0000110001110" => q_unbuf <= my_rom(398);
      when "0000110001111" => q_unbuf <= my_rom(399);
      when "0000110010000" => q_unbuf <= my_rom(400);
      when "0000110010001" => q_unbuf <= my_rom(401);
      when "0000110010010" => q_unbuf <= my_rom(402);
      when "0000110010011" => q_unbuf <= my_rom(403);
      when "0000110010100" => q_unbuf <= my_rom(404);
      when "0000110010101" => q_unbuf <= my_rom(405);
      when "0000110010110" => q_unbuf <= my_rom(406);
      when "0000110010111" => q_unbuf <= my_rom(407);
      when "0000110011000" => q_unbuf <= my_rom(408);
      when "0000110011001" => q_unbuf <= my_rom(409);
      when "0000110011010" => q_unbuf <= my_rom(410);
      when "0000110011011" => q_unbuf <= my_rom(411);
      when "0000110011100" => q_unbuf <= my_rom(412);
      when "0000110011101" => q_unbuf <= my_rom(413);
      when "0000110011110" => q_unbuf <= my_rom(414);
      when "0000110011111" => q_unbuf <= my_rom(415);
      when "0000110100000" => q_unbuf <= my_rom(416);
      when "0000110100001" => q_unbuf <= my_rom(417);
      when "0000110100010" => q_unbuf <= my_rom(418);
      when "0000110100011" => q_unbuf <= my_rom(419);
      when "0000110100100" => q_unbuf <= my_rom(420);
      when "0000110100101" => q_unbuf <= my_rom(421);
      when "0000110100110" => q_unbuf <= my_rom(422);
      when "0000110100111" => q_unbuf <= my_rom(423);
      when "0000110101000" => q_unbuf <= my_rom(424);
      when "0000110101001" => q_unbuf <= my_rom(425);
      when "0000110101010" => q_unbuf <= my_rom(426);
      when "0000110101011" => q_unbuf <= my_rom(427);
      when "0000110101100" => q_unbuf <= my_rom(428);
      when "0000110101101" => q_unbuf <= my_rom(429);
      when "0000110101110" => q_unbuf <= my_rom(430);
      when "0000110101111" => q_unbuf <= my_rom(431);
      when "0000110110000" => q_unbuf <= my_rom(432);
      when "0000110110001" => q_unbuf <= my_rom(433);
      when "0000110110010" => q_unbuf <= my_rom(434);
      when "0000110110011" => q_unbuf <= my_rom(435);
      when "0000110110100" => q_unbuf <= my_rom(436);
      when "0000110110101" => q_unbuf <= my_rom(437);
      when "0000110110110" => q_unbuf <= my_rom(438);
      when "0000110110111" => q_unbuf <= my_rom(439);
      when "0000110111000" => q_unbuf <= my_rom(440);
      when "0000110111001" => q_unbuf <= my_rom(441);
      when "0000110111010" => q_unbuf <= my_rom(442);
      when "0000110111011" => q_unbuf <= my_rom(443);
      when "0000110111100" => q_unbuf <= my_rom(444);
      when "0000110111101" => q_unbuf <= my_rom(445);
      when "0000110111110" => q_unbuf <= my_rom(446);
      when "0000110111111" => q_unbuf <= my_rom(447);
      when "0000111000000" => q_unbuf <= my_rom(448);
      when "0000111000001" => q_unbuf <= my_rom(449);
      when "0000111000010" => q_unbuf <= my_rom(450);
      when "0000111000011" => q_unbuf <= my_rom(451);
      when "0000111000100" => q_unbuf <= my_rom(452);
      when "0000111000101" => q_unbuf <= my_rom(453);
      when "0000111000110" => q_unbuf <= my_rom(454);
      when "0000111000111" => q_unbuf <= my_rom(455);
      when "0000111001000" => q_unbuf <= my_rom(456);
      when "0000111001001" => q_unbuf <= my_rom(457);
      when "0000111001010" => q_unbuf <= my_rom(458);
      when "0000111001011" => q_unbuf <= my_rom(459);
      when "0000111001100" => q_unbuf <= my_rom(460);
      when "0000111001101" => q_unbuf <= my_rom(461);
      when "0000111001110" => q_unbuf <= my_rom(462);
      when "0000111001111" => q_unbuf <= my_rom(463);
      when "0000111010000" => q_unbuf <= my_rom(464);
      when "0000111010001" => q_unbuf <= my_rom(465);
      when "0000111010010" => q_unbuf <= my_rom(466);
      when "0000111010011" => q_unbuf <= my_rom(467);
      when "0000111010100" => q_unbuf <= my_rom(468);
      when "0000111010101" => q_unbuf <= my_rom(469);
      when "0000111010110" => q_unbuf <= my_rom(470);
      when "0000111010111" => q_unbuf <= my_rom(471);
      when "0000111011000" => q_unbuf <= my_rom(472);
      when "0000111011001" => q_unbuf <= my_rom(473);
      when "0000111011010" => q_unbuf <= my_rom(474);
      when "0000111011011" => q_unbuf <= my_rom(475);
      when "0000111011100" => q_unbuf <= my_rom(476);
      when "0000111011101" => q_unbuf <= my_rom(477);
      when "0000111011110" => q_unbuf <= my_rom(478);
      when "0000111011111" => q_unbuf <= my_rom(479);
      when "0000111100000" => q_unbuf <= my_rom(480);
      when "0000111100001" => q_unbuf <= my_rom(481);
      when "0000111100010" => q_unbuf <= my_rom(482);
      when "0000111100011" => q_unbuf <= my_rom(483);
      when "0000111100100" => q_unbuf <= my_rom(484);
      when "0000111100101" => q_unbuf <= my_rom(485);
      when "0000111100110" => q_unbuf <= my_rom(486);
      when "0000111100111" => q_unbuf <= my_rom(487);
      when "0000111101000" => q_unbuf <= my_rom(488);
      when "0000111101001" => q_unbuf <= my_rom(489);
      when "0000111101010" => q_unbuf <= my_rom(490);
      when "0000111101011" => q_unbuf <= my_rom(491);
      when "0000111101100" => q_unbuf <= my_rom(492);
      when "0000111101101" => q_unbuf <= my_rom(493);
      when "0000111101110" => q_unbuf <= my_rom(494);
      when "0000111101111" => q_unbuf <= my_rom(495);
      when "0000111110000" => q_unbuf <= my_rom(496);
      when "0000111110001" => q_unbuf <= my_rom(497);
      when "0000111110010" => q_unbuf <= my_rom(498);
      when "0000111110011" => q_unbuf <= my_rom(499);
      when "0000111110100" => q_unbuf <= my_rom(500);
      when "0000111110101" => q_unbuf <= my_rom(501);
      when "0000111110110" => q_unbuf <= my_rom(502);
      when "0000111110111" => q_unbuf <= my_rom(503);
      when "0000111111000" => q_unbuf <= my_rom(504);
      when "0000111111001" => q_unbuf <= my_rom(505);
      when "0000111111010" => q_unbuf <= my_rom(506);
      when "0000111111011" => q_unbuf <= my_rom(507);
      when "0000111111100" => q_unbuf <= my_rom(508);
      when "0000111111101" => q_unbuf <= my_rom(509);
      when "0000111111110" => q_unbuf <= my_rom(510);
      when "0000111111111" => q_unbuf <= my_rom(511);
      when "0001000000000" => q_unbuf <= my_rom(512);
      when "0001000000001" => q_unbuf <= my_rom(513);
      when "0001000000010" => q_unbuf <= my_rom(514);
      when "0001000000011" => q_unbuf <= my_rom(515);
      when "0001000000100" => q_unbuf <= my_rom(516);
      when "0001000000101" => q_unbuf <= my_rom(517);
      when "0001000000110" => q_unbuf <= my_rom(518);
      when "0001000000111" => q_unbuf <= my_rom(519);
      when "0001000001000" => q_unbuf <= my_rom(520);
      when "0001000001001" => q_unbuf <= my_rom(521);
      when "0001000001010" => q_unbuf <= my_rom(522);
      when "0001000001011" => q_unbuf <= my_rom(523);
      when "0001000001100" => q_unbuf <= my_rom(524);
      when "0001000001101" => q_unbuf <= my_rom(525);
      when "0001000001110" => q_unbuf <= my_rom(526);
      when "0001000001111" => q_unbuf <= my_rom(527);
      when "0001000010000" => q_unbuf <= my_rom(528);
      when "0001000010001" => q_unbuf <= my_rom(529);
      when "0001000010010" => q_unbuf <= my_rom(530);
      when "0001000010011" => q_unbuf <= my_rom(531);
      when "0001000010100" => q_unbuf <= my_rom(532);
      when "0001000010101" => q_unbuf <= my_rom(533);
      when "0001000010110" => q_unbuf <= my_rom(534);
      when "0001000010111" => q_unbuf <= my_rom(535);
      when "0001000011000" => q_unbuf <= my_rom(536);
      when "0001000011001" => q_unbuf <= my_rom(537);
      when "0001000011010" => q_unbuf <= my_rom(538);
      when "0001000011011" => q_unbuf <= my_rom(539);
      when "0001000011100" => q_unbuf <= my_rom(540);
      when "0001000011101" => q_unbuf <= my_rom(541);
      when "0001000011110" => q_unbuf <= my_rom(542);
      when "0001000011111" => q_unbuf <= my_rom(543);
      when "0001000100000" => q_unbuf <= my_rom(544);
      when "0001000100001" => q_unbuf <= my_rom(545);
      when "0001000100010" => q_unbuf <= my_rom(546);
      when "0001000100011" => q_unbuf <= my_rom(547);
      when "0001000100100" => q_unbuf <= my_rom(548);
      when "0001000100101" => q_unbuf <= my_rom(549);
      when "0001000100110" => q_unbuf <= my_rom(550);
      when "0001000100111" => q_unbuf <= my_rom(551);
      when "0001000101000" => q_unbuf <= my_rom(552);
      when "0001000101001" => q_unbuf <= my_rom(553);
      when "0001000101010" => q_unbuf <= my_rom(554);
      when "0001000101011" => q_unbuf <= my_rom(555);
      when "0001000101100" => q_unbuf <= my_rom(556);
      when "0001000101101" => q_unbuf <= my_rom(557);
      when "0001000101110" => q_unbuf <= my_rom(558);
      when "0001000101111" => q_unbuf <= my_rom(559);
      when "0001000110000" => q_unbuf <= my_rom(560);
      when "0001000110001" => q_unbuf <= my_rom(561);
      when "0001000110010" => q_unbuf <= my_rom(562);
      when "0001000110011" => q_unbuf <= my_rom(563);
      when "0001000110100" => q_unbuf <= my_rom(564);
      when "0001000110101" => q_unbuf <= my_rom(565);
      when "0001000110110" => q_unbuf <= my_rom(566);
      when "0001000110111" => q_unbuf <= my_rom(567);
      when "0001000111000" => q_unbuf <= my_rom(568);
      when "0001000111001" => q_unbuf <= my_rom(569);
      when "0001000111010" => q_unbuf <= my_rom(570);
      when "0001000111011" => q_unbuf <= my_rom(571);
      when "0001000111100" => q_unbuf <= my_rom(572);
      when "0001000111101" => q_unbuf <= my_rom(573);
      when "0001000111110" => q_unbuf <= my_rom(574);
      when "0001000111111" => q_unbuf <= my_rom(575);
      when "0001001000000" => q_unbuf <= my_rom(576);
      when "0001001000001" => q_unbuf <= my_rom(577);
      when "0001001000010" => q_unbuf <= my_rom(578);
      when "0001001000011" => q_unbuf <= my_rom(579);
      when "0001001000100" => q_unbuf <= my_rom(580);
      when "0001001000101" => q_unbuf <= my_rom(581);
      when "0001001000110" => q_unbuf <= my_rom(582);
      when "0001001000111" => q_unbuf <= my_rom(583);
      when "0001001001000" => q_unbuf <= my_rom(584);
      when "0001001001001" => q_unbuf <= my_rom(585);
      when "0001001001010" => q_unbuf <= my_rom(586);
      when "0001001001011" => q_unbuf <= my_rom(587);
      when "0001001001100" => q_unbuf <= my_rom(588);
      when "0001001001101" => q_unbuf <= my_rom(589);
      when "0001001001110" => q_unbuf <= my_rom(590);
      when "0001001001111" => q_unbuf <= my_rom(591);
      when "0001001010000" => q_unbuf <= my_rom(592);
      when "0001001010001" => q_unbuf <= my_rom(593);
      when "0001001010010" => q_unbuf <= my_rom(594);
      when "0001001010011" => q_unbuf <= my_rom(595);
      when "0001001010100" => q_unbuf <= my_rom(596);
      when "0001001010101" => q_unbuf <= my_rom(597);
      when "0001001010110" => q_unbuf <= my_rom(598);
      when "0001001010111" => q_unbuf <= my_rom(599);
      when "0001001011000" => q_unbuf <= my_rom(600);
      when "0001001011001" => q_unbuf <= my_rom(601);
      when "0001001011010" => q_unbuf <= my_rom(602);
      when "0001001011011" => q_unbuf <= my_rom(603);
      when "0001001011100" => q_unbuf <= my_rom(604);
      when "0001001011101" => q_unbuf <= my_rom(605);
      when "0001001011110" => q_unbuf <= my_rom(606);
      when "0001001011111" => q_unbuf <= my_rom(607);
      when "0001001100000" => q_unbuf <= my_rom(608);
      when "0001001100001" => q_unbuf <= my_rom(609);
      when "0001001100010" => q_unbuf <= my_rom(610);
      when "0001001100011" => q_unbuf <= my_rom(611);
      when "0001001100100" => q_unbuf <= my_rom(612);
      when "0001001100101" => q_unbuf <= my_rom(613);
      when "0001001100110" => q_unbuf <= my_rom(614);
      when "0001001100111" => q_unbuf <= my_rom(615);
      when "0001001101000" => q_unbuf <= my_rom(616);
      when "0001001101001" => q_unbuf <= my_rom(617);
      when "0001001101010" => q_unbuf <= my_rom(618);
      when "0001001101011" => q_unbuf <= my_rom(619);
      when "0001001101100" => q_unbuf <= my_rom(620);
      when "0001001101101" => q_unbuf <= my_rom(621);
      when "0001001101110" => q_unbuf <= my_rom(622);
      when "0001001101111" => q_unbuf <= my_rom(623);
      when "0001001110000" => q_unbuf <= my_rom(624);
      when "0001001110001" => q_unbuf <= my_rom(625);
      when "0001001110010" => q_unbuf <= my_rom(626);
      when "0001001110011" => q_unbuf <= my_rom(627);
      when "0001001110100" => q_unbuf <= my_rom(628);
      when "0001001110101" => q_unbuf <= my_rom(629);
      when "0001001110110" => q_unbuf <= my_rom(630);
      when "0001001110111" => q_unbuf <= my_rom(631);
      when "0001001111000" => q_unbuf <= my_rom(632);
      when "0001001111001" => q_unbuf <= my_rom(633);
      when "0001001111010" => q_unbuf <= my_rom(634);
      when "0001001111011" => q_unbuf <= my_rom(635);
      when "0001001111100" => q_unbuf <= my_rom(636);
      when "0001001111101" => q_unbuf <= my_rom(637);
      when "0001001111110" => q_unbuf <= my_rom(638);
      when "0001001111111" => q_unbuf <= my_rom(639);
      when "0001010000000" => q_unbuf <= my_rom(640);
      when "0001010000001" => q_unbuf <= my_rom(641);
      when "0001010000010" => q_unbuf <= my_rom(642);
      when "0001010000011" => q_unbuf <= my_rom(643);
      when "0001010000100" => q_unbuf <= my_rom(644);
      when "0001010000101" => q_unbuf <= my_rom(645);
      when "0001010000110" => q_unbuf <= my_rom(646);
      when "0001010000111" => q_unbuf <= my_rom(647);
      when "0001010001000" => q_unbuf <= my_rom(648);
      when "0001010001001" => q_unbuf <= my_rom(649);
      when "0001010001010" => q_unbuf <= my_rom(650);
      when "0001010001011" => q_unbuf <= my_rom(651);
      when "0001010001100" => q_unbuf <= my_rom(652);
      when "0001010001101" => q_unbuf <= my_rom(653);
      when "0001010001110" => q_unbuf <= my_rom(654);
      when "0001010001111" => q_unbuf <= my_rom(655);
      when "0001010010000" => q_unbuf <= my_rom(656);
      when "0001010010001" => q_unbuf <= my_rom(657);
      when "0001010010010" => q_unbuf <= my_rom(658);
      when "0001010010011" => q_unbuf <= my_rom(659);
      when "0001010010100" => q_unbuf <= my_rom(660);
      when "0001010010101" => q_unbuf <= my_rom(661);
      when "0001010010110" => q_unbuf <= my_rom(662);
      when "0001010010111" => q_unbuf <= my_rom(663);
      when "0001010011000" => q_unbuf <= my_rom(664);
      when "0001010011001" => q_unbuf <= my_rom(665);
      when "0001010011010" => q_unbuf <= my_rom(666);
      when "0001010011011" => q_unbuf <= my_rom(667);
      when "0001010011100" => q_unbuf <= my_rom(668);
      when "0001010011101" => q_unbuf <= my_rom(669);
      when "0001010011110" => q_unbuf <= my_rom(670);
      when "0001010011111" => q_unbuf <= my_rom(671);
      when "0001010100000" => q_unbuf <= my_rom(672);
      when "0001010100001" => q_unbuf <= my_rom(673);
      when "0001010100010" => q_unbuf <= my_rom(674);
      when "0001010100011" => q_unbuf <= my_rom(675);
      when "0001010100100" => q_unbuf <= my_rom(676);
      when "0001010100101" => q_unbuf <= my_rom(677);
      when "0001010100110" => q_unbuf <= my_rom(678);
      when "0001010100111" => q_unbuf <= my_rom(679);
      when "0001010101000" => q_unbuf <= my_rom(680);
      when "0001010101001" => q_unbuf <= my_rom(681);
      when "0001010101010" => q_unbuf <= my_rom(682);
      when "0001010101011" => q_unbuf <= my_rom(683);
      when "0001010101100" => q_unbuf <= my_rom(684);
      when "0001010101101" => q_unbuf <= my_rom(685);
      when "0001010101110" => q_unbuf <= my_rom(686);
      when "0001010101111" => q_unbuf <= my_rom(687);
      when "0001010110000" => q_unbuf <= my_rom(688);
      when "0001010110001" => q_unbuf <= my_rom(689);
      when "0001010110010" => q_unbuf <= my_rom(690);
      when "0001010110011" => q_unbuf <= my_rom(691);
      when "0001010110100" => q_unbuf <= my_rom(692);
      when "0001010110101" => q_unbuf <= my_rom(693);
      when "0001010110110" => q_unbuf <= my_rom(694);
      when "0001010110111" => q_unbuf <= my_rom(695);
      when "0001010111000" => q_unbuf <= my_rom(696);
      when "0001010111001" => q_unbuf <= my_rom(697);
      when "0001010111010" => q_unbuf <= my_rom(698);
      when "0001010111011" => q_unbuf <= my_rom(699);
      when "0001010111100" => q_unbuf <= my_rom(700);
      when "0001010111101" => q_unbuf <= my_rom(701);
      when "0001010111110" => q_unbuf <= my_rom(702);
      when "0001010111111" => q_unbuf <= my_rom(703);
      when "0001011000000" => q_unbuf <= my_rom(704);
      when "0001011000001" => q_unbuf <= my_rom(705);
      when "0001011000010" => q_unbuf <= my_rom(706);
      when "0001011000011" => q_unbuf <= my_rom(707);
      when "0001011000100" => q_unbuf <= my_rom(708);
      when "0001011000101" => q_unbuf <= my_rom(709);
      when "0001011000110" => q_unbuf <= my_rom(710);
      when "0001011000111" => q_unbuf <= my_rom(711);
      when "0001011001000" => q_unbuf <= my_rom(712);
      when "0001011001001" => q_unbuf <= my_rom(713);
      when "0001011001010" => q_unbuf <= my_rom(714);
      when "0001011001011" => q_unbuf <= my_rom(715);
      when "0001011001100" => q_unbuf <= my_rom(716);
      when "0001011001101" => q_unbuf <= my_rom(717);
      when "0001011001110" => q_unbuf <= my_rom(718);
      when "0001011001111" => q_unbuf <= my_rom(719);
      when "0001011010000" => q_unbuf <= my_rom(720);
      when "0001011010001" => q_unbuf <= my_rom(721);
      when "0001011010010" => q_unbuf <= my_rom(722);
      when "0001011010011" => q_unbuf <= my_rom(723);
      when "0001011010100" => q_unbuf <= my_rom(724);
      when "0001011010101" => q_unbuf <= my_rom(725);
      when "0001011010110" => q_unbuf <= my_rom(726);
      when "0001011010111" => q_unbuf <= my_rom(727);
      when "0001011011000" => q_unbuf <= my_rom(728);
      when "0001011011001" => q_unbuf <= my_rom(729);
      when "0001011011010" => q_unbuf <= my_rom(730);
      when "0001011011011" => q_unbuf <= my_rom(731);
      when "0001011011100" => q_unbuf <= my_rom(732);
      when "0001011011101" => q_unbuf <= my_rom(733);
      when "0001011011110" => q_unbuf <= my_rom(734);
      when "0001011011111" => q_unbuf <= my_rom(735);
      when "0001011100000" => q_unbuf <= my_rom(736);
      when "0001011100001" => q_unbuf <= my_rom(737);
      when "0001011100010" => q_unbuf <= my_rom(738);
      when "0001011100011" => q_unbuf <= my_rom(739);
      when "0001011100100" => q_unbuf <= my_rom(740);
      when "0001011100101" => q_unbuf <= my_rom(741);
      when "0001011100110" => q_unbuf <= my_rom(742);
      when "0001011100111" => q_unbuf <= my_rom(743);
      when "0001011101000" => q_unbuf <= my_rom(744);
      when "0001011101001" => q_unbuf <= my_rom(745);
      when "0001011101010" => q_unbuf <= my_rom(746);
      when "0001011101011" => q_unbuf <= my_rom(747);
      when "0001011101100" => q_unbuf <= my_rom(748);
      when "0001011101101" => q_unbuf <= my_rom(749);
      when "0001011101110" => q_unbuf <= my_rom(750);
      when "0001011101111" => q_unbuf <= my_rom(751);
      when "0001011110000" => q_unbuf <= my_rom(752);
      when "0001011110001" => q_unbuf <= my_rom(753);
      when "0001011110010" => q_unbuf <= my_rom(754);
      when "0001011110011" => q_unbuf <= my_rom(755);
      when "0001011110100" => q_unbuf <= my_rom(756);
      when "0001011110101" => q_unbuf <= my_rom(757);
      when "0001011110110" => q_unbuf <= my_rom(758);
      when "0001011110111" => q_unbuf <= my_rom(759);
      when "0001011111000" => q_unbuf <= my_rom(760);
      when "0001011111001" => q_unbuf <= my_rom(761);
      when "0001011111010" => q_unbuf <= my_rom(762);
      when "0001011111011" => q_unbuf <= my_rom(763);
      when "0001011111100" => q_unbuf <= my_rom(764);
      when "0001011111101" => q_unbuf <= my_rom(765);
      when "0001011111110" => q_unbuf <= my_rom(766);
      when "0001011111111" => q_unbuf <= my_rom(767);
      when "0001100000000" => q_unbuf <= my_rom(768);
      when "0001100000001" => q_unbuf <= my_rom(769);
      when "0001100000010" => q_unbuf <= my_rom(770);
      when "0001100000011" => q_unbuf <= my_rom(771);
      when "0001100000100" => q_unbuf <= my_rom(772);
      when "0001100000101" => q_unbuf <= my_rom(773);
      when "0001100000110" => q_unbuf <= my_rom(774);
      when "0001100000111" => q_unbuf <= my_rom(775);
      when "0001100001000" => q_unbuf <= my_rom(776);
      when "0001100001001" => q_unbuf <= my_rom(777);
      when "0001100001010" => q_unbuf <= my_rom(778);
      when "0001100001011" => q_unbuf <= my_rom(779);
      when "0001100001100" => q_unbuf <= my_rom(780);
      when "0001100001101" => q_unbuf <= my_rom(781);
      when "0001100001110" => q_unbuf <= my_rom(782);
      when "0001100001111" => q_unbuf <= my_rom(783);
      when "0001100010000" => q_unbuf <= my_rom(784);
      when "0001100010001" => q_unbuf <= my_rom(785);
      when "0001100010010" => q_unbuf <= my_rom(786);
      when "0001100010011" => q_unbuf <= my_rom(787);
      when "0001100010100" => q_unbuf <= my_rom(788);
      when "0001100010101" => q_unbuf <= my_rom(789);
      when "0001100010110" => q_unbuf <= my_rom(790);
      when "0001100010111" => q_unbuf <= my_rom(791);
      when "0001100011000" => q_unbuf <= my_rom(792);
      when "0001100011001" => q_unbuf <= my_rom(793);
      when "0001100011010" => q_unbuf <= my_rom(794);
      when "0001100011011" => q_unbuf <= my_rom(795);
      when "0001100011100" => q_unbuf <= my_rom(796);
      when "0001100011101" => q_unbuf <= my_rom(797);
      when "0001100011110" => q_unbuf <= my_rom(798);
      when "0001100011111" => q_unbuf <= my_rom(799);
      when "0001100100000" => q_unbuf <= my_rom(800);
      when "0001100100001" => q_unbuf <= my_rom(801);
      when "0001100100010" => q_unbuf <= my_rom(802);
      when "0001100100011" => q_unbuf <= my_rom(803);
      when "0001100100100" => q_unbuf <= my_rom(804);
      when "0001100100101" => q_unbuf <= my_rom(805);
      when "0001100100110" => q_unbuf <= my_rom(806);
      when "0001100100111" => q_unbuf <= my_rom(807);
      when "0001100101000" => q_unbuf <= my_rom(808);
      when "0001100101001" => q_unbuf <= my_rom(809);
      when "0001100101010" => q_unbuf <= my_rom(810);
      when "0001100101011" => q_unbuf <= my_rom(811);
      when "0001100101100" => q_unbuf <= my_rom(812);
      when "0001100101101" => q_unbuf <= my_rom(813);
      when "0001100101110" => q_unbuf <= my_rom(814);
      when "0001100101111" => q_unbuf <= my_rom(815);
      when "0001100110000" => q_unbuf <= my_rom(816);
      when "0001100110001" => q_unbuf <= my_rom(817);
      when "0001100110010" => q_unbuf <= my_rom(818);
      when "0001100110011" => q_unbuf <= my_rom(819);
      when "0001100110100" => q_unbuf <= my_rom(820);
      when "0001100110101" => q_unbuf <= my_rom(821);
      when "0001100110110" => q_unbuf <= my_rom(822);
      when "0001100110111" => q_unbuf <= my_rom(823);
      when "0001100111000" => q_unbuf <= my_rom(824);
      when "0001100111001" => q_unbuf <= my_rom(825);
      when "0001100111010" => q_unbuf <= my_rom(826);
      when "0001100111011" => q_unbuf <= my_rom(827);
      when "0001100111100" => q_unbuf <= my_rom(828);
      when "0001100111101" => q_unbuf <= my_rom(829);
      when "0001100111110" => q_unbuf <= my_rom(830);
      when "0001100111111" => q_unbuf <= my_rom(831);
      when "0001101000000" => q_unbuf <= my_rom(832);
      when "0001101000001" => q_unbuf <= my_rom(833);
      when "0001101000010" => q_unbuf <= my_rom(834);
      when "0001101000011" => q_unbuf <= my_rom(835);
      when "0001101000100" => q_unbuf <= my_rom(836);
      when "0001101000101" => q_unbuf <= my_rom(837);
      when "0001101000110" => q_unbuf <= my_rom(838);
      when "0001101000111" => q_unbuf <= my_rom(839);
      when "0001101001000" => q_unbuf <= my_rom(840);
      when "0001101001001" => q_unbuf <= my_rom(841);
      when "0001101001010" => q_unbuf <= my_rom(842);
      when "0001101001011" => q_unbuf <= my_rom(843);
      when "0001101001100" => q_unbuf <= my_rom(844);
      when "0001101001101" => q_unbuf <= my_rom(845);
      when "0001101001110" => q_unbuf <= my_rom(846);
      when "0001101001111" => q_unbuf <= my_rom(847);
      when "0001101010000" => q_unbuf <= my_rom(848);
      when "0001101010001" => q_unbuf <= my_rom(849);
      when "0001101010010" => q_unbuf <= my_rom(850);
      when "0001101010011" => q_unbuf <= my_rom(851);
      when "0001101010100" => q_unbuf <= my_rom(852);
      when "0001101010101" => q_unbuf <= my_rom(853);
      when "0001101010110" => q_unbuf <= my_rom(854);
      when "0001101010111" => q_unbuf <= my_rom(855);
      when "0001101011000" => q_unbuf <= my_rom(856);
      when "0001101011001" => q_unbuf <= my_rom(857);
      when "0001101011010" => q_unbuf <= my_rom(858);
      when "0001101011011" => q_unbuf <= my_rom(859);
      when "0001101011100" => q_unbuf <= my_rom(860);
      when "0001101011101" => q_unbuf <= my_rom(861);
      when "0001101011110" => q_unbuf <= my_rom(862);
      when "0001101011111" => q_unbuf <= my_rom(863);
      when "0001101100000" => q_unbuf <= my_rom(864);
      when "0001101100001" => q_unbuf <= my_rom(865);
      when "0001101100010" => q_unbuf <= my_rom(866);
      when "0001101100011" => q_unbuf <= my_rom(867);
      when "0001101100100" => q_unbuf <= my_rom(868);
      when "0001101100101" => q_unbuf <= my_rom(869);
      when "0001101100110" => q_unbuf <= my_rom(870);
      when "0001101100111" => q_unbuf <= my_rom(871);
      when "0001101101000" => q_unbuf <= my_rom(872);
      when "0001101101001" => q_unbuf <= my_rom(873);
      when "0001101101010" => q_unbuf <= my_rom(874);
      when "0001101101011" => q_unbuf <= my_rom(875);
      when "0001101101100" => q_unbuf <= my_rom(876);
      when "0001101101101" => q_unbuf <= my_rom(877);
      when "0001101101110" => q_unbuf <= my_rom(878);
      when "0001101101111" => q_unbuf <= my_rom(879);
      when "0001101110000" => q_unbuf <= my_rom(880);
      when "0001101110001" => q_unbuf <= my_rom(881);
      when "0001101110010" => q_unbuf <= my_rom(882);
      when "0001101110011" => q_unbuf <= my_rom(883);
      when "0001101110100" => q_unbuf <= my_rom(884);
      when "0001101110101" => q_unbuf <= my_rom(885);
      when "0001101110110" => q_unbuf <= my_rom(886);
      when "0001101110111" => q_unbuf <= my_rom(887);
      when "0001101111000" => q_unbuf <= my_rom(888);
      when "0001101111001" => q_unbuf <= my_rom(889);
      when "0001101111010" => q_unbuf <= my_rom(890);
      when "0001101111011" => q_unbuf <= my_rom(891);
      when "0001101111100" => q_unbuf <= my_rom(892);
      when "0001101111101" => q_unbuf <= my_rom(893);
      when "0001101111110" => q_unbuf <= my_rom(894);
      when "0001101111111" => q_unbuf <= my_rom(895);
      when "0001110000000" => q_unbuf <= my_rom(896);
      when "0001110000001" => q_unbuf <= my_rom(897);
      when "0001110000010" => q_unbuf <= my_rom(898);
      when "0001110000011" => q_unbuf <= my_rom(899);
      when "0001110000100" => q_unbuf <= my_rom(900);
      when "0001110000101" => q_unbuf <= my_rom(901);
      when "0001110000110" => q_unbuf <= my_rom(902);
      when "0001110000111" => q_unbuf <= my_rom(903);
      when "0001110001000" => q_unbuf <= my_rom(904);
      when "0001110001001" => q_unbuf <= my_rom(905);
      when "0001110001010" => q_unbuf <= my_rom(906);
      when "0001110001011" => q_unbuf <= my_rom(907);
      when "0001110001100" => q_unbuf <= my_rom(908);
      when "0001110001101" => q_unbuf <= my_rom(909);
      when "0001110001110" => q_unbuf <= my_rom(910);
      when "0001110001111" => q_unbuf <= my_rom(911);
      when "0001110010000" => q_unbuf <= my_rom(912);
      when "0001110010001" => q_unbuf <= my_rom(913);
      when "0001110010010" => q_unbuf <= my_rom(914);
      when "0001110010011" => q_unbuf <= my_rom(915);
      when "0001110010100" => q_unbuf <= my_rom(916);
      when "0001110010101" => q_unbuf <= my_rom(917);
      when "0001110010110" => q_unbuf <= my_rom(918);
      when "0001110010111" => q_unbuf <= my_rom(919);
      when "0001110011000" => q_unbuf <= my_rom(920);
      when "0001110011001" => q_unbuf <= my_rom(921);
      when "0001110011010" => q_unbuf <= my_rom(922);
      when "0001110011011" => q_unbuf <= my_rom(923);
      when "0001110011100" => q_unbuf <= my_rom(924);
      when "0001110011101" => q_unbuf <= my_rom(925);
      when "0001110011110" => q_unbuf <= my_rom(926);
      when "0001110011111" => q_unbuf <= my_rom(927);
      when "0001110100000" => q_unbuf <= my_rom(928);
      when "0001110100001" => q_unbuf <= my_rom(929);
      when "0001110100010" => q_unbuf <= my_rom(930);
      when "0001110100011" => q_unbuf <= my_rom(931);
      when "0001110100100" => q_unbuf <= my_rom(932);
      when "0001110100101" => q_unbuf <= my_rom(933);
      when "0001110100110" => q_unbuf <= my_rom(934);
      when "0001110100111" => q_unbuf <= my_rom(935);
      when "0001110101000" => q_unbuf <= my_rom(936);
      when "0001110101001" => q_unbuf <= my_rom(937);
      when "0001110101010" => q_unbuf <= my_rom(938);
      when "0001110101011" => q_unbuf <= my_rom(939);
      when "0001110101100" => q_unbuf <= my_rom(940);
      when "0001110101101" => q_unbuf <= my_rom(941);
      when "0001110101110" => q_unbuf <= my_rom(942);
      when "0001110101111" => q_unbuf <= my_rom(943);
      when "0001110110000" => q_unbuf <= my_rom(944);
      when "0001110110001" => q_unbuf <= my_rom(945);
      when "0001110110010" => q_unbuf <= my_rom(946);
      when "0001110110011" => q_unbuf <= my_rom(947);
      when "0001110110100" => q_unbuf <= my_rom(948);
      when "0001110110101" => q_unbuf <= my_rom(949);
      when "0001110110110" => q_unbuf <= my_rom(950);
      when "0001110110111" => q_unbuf <= my_rom(951);
      when "0001110111000" => q_unbuf <= my_rom(952);
      when "0001110111001" => q_unbuf <= my_rom(953);
      when "0001110111010" => q_unbuf <= my_rom(954);
      when "0001110111011" => q_unbuf <= my_rom(955);
      when "0001110111100" => q_unbuf <= my_rom(956);
      when "0001110111101" => q_unbuf <= my_rom(957);
      when "0001110111110" => q_unbuf <= my_rom(958);
      when "0001110111111" => q_unbuf <= my_rom(959);
      when "0001111000000" => q_unbuf <= my_rom(960);
      when "0001111000001" => q_unbuf <= my_rom(961);
      when "0001111000010" => q_unbuf <= my_rom(962);
      when "0001111000011" => q_unbuf <= my_rom(963);
      when "0001111000100" => q_unbuf <= my_rom(964);
      when "0001111000101" => q_unbuf <= my_rom(965);
      when "0001111000110" => q_unbuf <= my_rom(966);
      when "0001111000111" => q_unbuf <= my_rom(967);
      when "0001111001000" => q_unbuf <= my_rom(968);
      when "0001111001001" => q_unbuf <= my_rom(969);
      when "0001111001010" => q_unbuf <= my_rom(970);
      when "0001111001011" => q_unbuf <= my_rom(971);
      when "0001111001100" => q_unbuf <= my_rom(972);
      when "0001111001101" => q_unbuf <= my_rom(973);
      when "0001111001110" => q_unbuf <= my_rom(974);
      when "0001111001111" => q_unbuf <= my_rom(975);
      when "0001111010000" => q_unbuf <= my_rom(976);
      when "0001111010001" => q_unbuf <= my_rom(977);
      when "0001111010010" => q_unbuf <= my_rom(978);
      when "0001111010011" => q_unbuf <= my_rom(979);
      when "0001111010100" => q_unbuf <= my_rom(980);
      when "0001111010101" => q_unbuf <= my_rom(981);
      when "0001111010110" => q_unbuf <= my_rom(982);
      when "0001111010111" => q_unbuf <= my_rom(983);
      when "0001111011000" => q_unbuf <= my_rom(984);
      when "0001111011001" => q_unbuf <= my_rom(985);
      when "0001111011010" => q_unbuf <= my_rom(986);
      when "0001111011011" => q_unbuf <= my_rom(987);
      when "0001111011100" => q_unbuf <= my_rom(988);
      when "0001111011101" => q_unbuf <= my_rom(989);
      when "0001111011110" => q_unbuf <= my_rom(990);
      when "0001111011111" => q_unbuf <= my_rom(991);
      when "0001111100000" => q_unbuf <= my_rom(992);
      when "0001111100001" => q_unbuf <= my_rom(993);
      when "0001111100010" => q_unbuf <= my_rom(994);
      when "0001111100011" => q_unbuf <= my_rom(995);
      when "0001111100100" => q_unbuf <= my_rom(996);
      when "0001111100101" => q_unbuf <= my_rom(997);
      when "0001111100110" => q_unbuf <= my_rom(998);
      when "0001111100111" => q_unbuf <= my_rom(999);
      when "0001111101000" => q_unbuf <= my_rom(1000);
      when "0001111101001" => q_unbuf <= my_rom(1001);
      when "0001111101010" => q_unbuf <= my_rom(1002);
      when "0001111101011" => q_unbuf <= my_rom(1003);
      when "0001111101100" => q_unbuf <= my_rom(1004);
      when "0001111101101" => q_unbuf <= my_rom(1005);
      when "0001111101110" => q_unbuf <= my_rom(1006);
      when "0001111101111" => q_unbuf <= my_rom(1007);
      when "0001111110000" => q_unbuf <= my_rom(1008);
      when "0001111110001" => q_unbuf <= my_rom(1009);
      when "0001111110010" => q_unbuf <= my_rom(1010);
      when "0001111110011" => q_unbuf <= my_rom(1011);
      when "0001111110100" => q_unbuf <= my_rom(1012);
      when "0001111110101" => q_unbuf <= my_rom(1013);
      when "0001111110110" => q_unbuf <= my_rom(1014);
      when "0001111110111" => q_unbuf <= my_rom(1015);
      when "0001111111000" => q_unbuf <= my_rom(1016);
      when "0001111111001" => q_unbuf <= my_rom(1017);
      when "0001111111010" => q_unbuf <= my_rom(1018);
      when "0001111111011" => q_unbuf <= my_rom(1019);
      when "0001111111100" => q_unbuf <= my_rom(1020);
      when "0001111111101" => q_unbuf <= my_rom(1021);
      when "0001111111110" => q_unbuf <= my_rom(1022);
      when "0001111111111" => q_unbuf <= my_rom(1023);
      when "0010000000000" => q_unbuf <= my_rom(1024);
      when "0010000000001" => q_unbuf <= my_rom(1025);
      when "0010000000010" => q_unbuf <= my_rom(1026);
      when "0010000000011" => q_unbuf <= my_rom(1027);
      when "0010000000100" => q_unbuf <= my_rom(1028);
      when "0010000000101" => q_unbuf <= my_rom(1029);
      when "0010000000110" => q_unbuf <= my_rom(1030);
      when "0010000000111" => q_unbuf <= my_rom(1031);
      when "0010000001000" => q_unbuf <= my_rom(1032);
      when "0010000001001" => q_unbuf <= my_rom(1033);
      when "0010000001010" => q_unbuf <= my_rom(1034);
      when "0010000001011" => q_unbuf <= my_rom(1035);
      when "0010000001100" => q_unbuf <= my_rom(1036);
      when "0010000001101" => q_unbuf <= my_rom(1037);
      when "0010000001110" => q_unbuf <= my_rom(1038);
      when "0010000001111" => q_unbuf <= my_rom(1039);
      when "0010000010000" => q_unbuf <= my_rom(1040);
      when "0010000010001" => q_unbuf <= my_rom(1041);
      when "0010000010010" => q_unbuf <= my_rom(1042);
      when "0010000010011" => q_unbuf <= my_rom(1043);
      when "0010000010100" => q_unbuf <= my_rom(1044);
      when "0010000010101" => q_unbuf <= my_rom(1045);
      when "0010000010110" => q_unbuf <= my_rom(1046);
      when "0010000010111" => q_unbuf <= my_rom(1047);
      when "0010000011000" => q_unbuf <= my_rom(1048);
      when "0010000011001" => q_unbuf <= my_rom(1049);
      when "0010000011010" => q_unbuf <= my_rom(1050);
      when "0010000011011" => q_unbuf <= my_rom(1051);
      when "0010000011100" => q_unbuf <= my_rom(1052);
      when "0010000011101" => q_unbuf <= my_rom(1053);
      when "0010000011110" => q_unbuf <= my_rom(1054);
      when "0010000011111" => q_unbuf <= my_rom(1055);
      when "0010000100000" => q_unbuf <= my_rom(1056);
      when "0010000100001" => q_unbuf <= my_rom(1057);
      when "0010000100010" => q_unbuf <= my_rom(1058);
      when "0010000100011" => q_unbuf <= my_rom(1059);
      when "0010000100100" => q_unbuf <= my_rom(1060);
      when "0010000100101" => q_unbuf <= my_rom(1061);
      when "0010000100110" => q_unbuf <= my_rom(1062);
      when "0010000100111" => q_unbuf <= my_rom(1063);
      when "0010000101000" => q_unbuf <= my_rom(1064);
      when "0010000101001" => q_unbuf <= my_rom(1065);
      when "0010000101010" => q_unbuf <= my_rom(1066);
      when "0010000101011" => q_unbuf <= my_rom(1067);
      when "0010000101100" => q_unbuf <= my_rom(1068);
      when "0010000101101" => q_unbuf <= my_rom(1069);
      when "0010000101110" => q_unbuf <= my_rom(1070);
      when "0010000101111" => q_unbuf <= my_rom(1071);
      when "0010000110000" => q_unbuf <= my_rom(1072);
      when "0010000110001" => q_unbuf <= my_rom(1073);
      when "0010000110010" => q_unbuf <= my_rom(1074);
      when "0010000110011" => q_unbuf <= my_rom(1075);
      when "0010000110100" => q_unbuf <= my_rom(1076);
      when "0010000110101" => q_unbuf <= my_rom(1077);
      when "0010000110110" => q_unbuf <= my_rom(1078);
      when "0010000110111" => q_unbuf <= my_rom(1079);
      when "0010000111000" => q_unbuf <= my_rom(1080);
      when "0010000111001" => q_unbuf <= my_rom(1081);
      when "0010000111010" => q_unbuf <= my_rom(1082);
      when "0010000111011" => q_unbuf <= my_rom(1083);
      when "0010000111100" => q_unbuf <= my_rom(1084);
      when "0010000111101" => q_unbuf <= my_rom(1085);
      when "0010000111110" => q_unbuf <= my_rom(1086);
      when "0010000111111" => q_unbuf <= my_rom(1087);
      when "0010001000000" => q_unbuf <= my_rom(1088);
      when "0010001000001" => q_unbuf <= my_rom(1089);
      when "0010001000010" => q_unbuf <= my_rom(1090);
      when "0010001000011" => q_unbuf <= my_rom(1091);
      when "0010001000100" => q_unbuf <= my_rom(1092);
      when "0010001000101" => q_unbuf <= my_rom(1093);
      when "0010001000110" => q_unbuf <= my_rom(1094);
      when "0010001000111" => q_unbuf <= my_rom(1095);
      when "0010001001000" => q_unbuf <= my_rom(1096);
      when "0010001001001" => q_unbuf <= my_rom(1097);
      when "0010001001010" => q_unbuf <= my_rom(1098);
      when "0010001001011" => q_unbuf <= my_rom(1099);
      when "0010001001100" => q_unbuf <= my_rom(1100);
      when "0010001001101" => q_unbuf <= my_rom(1101);
      when "0010001001110" => q_unbuf <= my_rom(1102);
      when "0010001001111" => q_unbuf <= my_rom(1103);
      when "0010001010000" => q_unbuf <= my_rom(1104);
      when "0010001010001" => q_unbuf <= my_rom(1105);
      when "0010001010010" => q_unbuf <= my_rom(1106);
      when "0010001010011" => q_unbuf <= my_rom(1107);
      when "0010001010100" => q_unbuf <= my_rom(1108);
      when "0010001010101" => q_unbuf <= my_rom(1109);
      when "0010001010110" => q_unbuf <= my_rom(1110);
      when "0010001010111" => q_unbuf <= my_rom(1111);
      when "0010001011000" => q_unbuf <= my_rom(1112);
      when "0010001011001" => q_unbuf <= my_rom(1113);
      when "0010001011010" => q_unbuf <= my_rom(1114);
      when "0010001011011" => q_unbuf <= my_rom(1115);
      when "0010001011100" => q_unbuf <= my_rom(1116);
      when "0010001011101" => q_unbuf <= my_rom(1117);
      when "0010001011110" => q_unbuf <= my_rom(1118);
      when "0010001011111" => q_unbuf <= my_rom(1119);
      when "0010001100000" => q_unbuf <= my_rom(1120);
      when "0010001100001" => q_unbuf <= my_rom(1121);
      when "0010001100010" => q_unbuf <= my_rom(1122);
      when "0010001100011" => q_unbuf <= my_rom(1123);
      when "0010001100100" => q_unbuf <= my_rom(1124);
      when "0010001100101" => q_unbuf <= my_rom(1125);
      when "0010001100110" => q_unbuf <= my_rom(1126);
      when "0010001100111" => q_unbuf <= my_rom(1127);
      when "0010001101000" => q_unbuf <= my_rom(1128);
      when "0010001101001" => q_unbuf <= my_rom(1129);
      when "0010001101010" => q_unbuf <= my_rom(1130);
      when "0010001101011" => q_unbuf <= my_rom(1131);
      when "0010001101100" => q_unbuf <= my_rom(1132);
      when "0010001101101" => q_unbuf <= my_rom(1133);
      when "0010001101110" => q_unbuf <= my_rom(1134);
      when "0010001101111" => q_unbuf <= my_rom(1135);
      when "0010001110000" => q_unbuf <= my_rom(1136);
      when "0010001110001" => q_unbuf <= my_rom(1137);
      when "0010001110010" => q_unbuf <= my_rom(1138);
      when "0010001110011" => q_unbuf <= my_rom(1139);
      when "0010001110100" => q_unbuf <= my_rom(1140);
      when "0010001110101" => q_unbuf <= my_rom(1141);
      when "0010001110110" => q_unbuf <= my_rom(1142);
      when "0010001110111" => q_unbuf <= my_rom(1143);
      when "0010001111000" => q_unbuf <= my_rom(1144);
      when "0010001111001" => q_unbuf <= my_rom(1145);
      when "0010001111010" => q_unbuf <= my_rom(1146);
      when "0010001111011" => q_unbuf <= my_rom(1147);
      when "0010001111100" => q_unbuf <= my_rom(1148);
      when "0010001111101" => q_unbuf <= my_rom(1149);
      when "0010001111110" => q_unbuf <= my_rom(1150);
      when "0010001111111" => q_unbuf <= my_rom(1151);
      when "0010010000000" => q_unbuf <= my_rom(1152);
      when "0010010000001" => q_unbuf <= my_rom(1153);
      when "0010010000010" => q_unbuf <= my_rom(1154);
      when "0010010000011" => q_unbuf <= my_rom(1155);
      when "0010010000100" => q_unbuf <= my_rom(1156);
      when "0010010000101" => q_unbuf <= my_rom(1157);
      when "0010010000110" => q_unbuf <= my_rom(1158);
      when "0010010000111" => q_unbuf <= my_rom(1159);
      when "0010010001000" => q_unbuf <= my_rom(1160);
      when "0010010001001" => q_unbuf <= my_rom(1161);
      when "0010010001010" => q_unbuf <= my_rom(1162);
      when "0010010001011" => q_unbuf <= my_rom(1163);
      when "0010010001100" => q_unbuf <= my_rom(1164);
      when "0010010001101" => q_unbuf <= my_rom(1165);
      when "0010010001110" => q_unbuf <= my_rom(1166);
      when "0010010001111" => q_unbuf <= my_rom(1167);
      when "0010010010000" => q_unbuf <= my_rom(1168);
      when "0010010010001" => q_unbuf <= my_rom(1169);
      when "0010010010010" => q_unbuf <= my_rom(1170);
      when "0010010010011" => q_unbuf <= my_rom(1171);
      when "0010010010100" => q_unbuf <= my_rom(1172);
      when "0010010010101" => q_unbuf <= my_rom(1173);
      when "0010010010110" => q_unbuf <= my_rom(1174);
      when "0010010010111" => q_unbuf <= my_rom(1175);
      when "0010010011000" => q_unbuf <= my_rom(1176);
      when "0010010011001" => q_unbuf <= my_rom(1177);
      when "0010010011010" => q_unbuf <= my_rom(1178);
      when "0010010011011" => q_unbuf <= my_rom(1179);
      when "0010010011100" => q_unbuf <= my_rom(1180);
      when "0010010011101" => q_unbuf <= my_rom(1181);
      when "0010010011110" => q_unbuf <= my_rom(1182);
      when "0010010011111" => q_unbuf <= my_rom(1183);
      when "0010010100000" => q_unbuf <= my_rom(1184);
      when "0010010100001" => q_unbuf <= my_rom(1185);
      when "0010010100010" => q_unbuf <= my_rom(1186);
      when "0010010100011" => q_unbuf <= my_rom(1187);
      when "0010010100100" => q_unbuf <= my_rom(1188);
      when "0010010100101" => q_unbuf <= my_rom(1189);
      when "0010010100110" => q_unbuf <= my_rom(1190);
      when "0010010100111" => q_unbuf <= my_rom(1191);
      when "0010010101000" => q_unbuf <= my_rom(1192);
      when "0010010101001" => q_unbuf <= my_rom(1193);
      when "0010010101010" => q_unbuf <= my_rom(1194);
      when "0010010101011" => q_unbuf <= my_rom(1195);
      when "0010010101100" => q_unbuf <= my_rom(1196);
      when "0010010101101" => q_unbuf <= my_rom(1197);
      when "0010010101110" => q_unbuf <= my_rom(1198);
      when "0010010101111" => q_unbuf <= my_rom(1199);
      when "0010010110000" => q_unbuf <= my_rom(1200);
      when "0010010110001" => q_unbuf <= my_rom(1201);
      when "0010010110010" => q_unbuf <= my_rom(1202);
      when "0010010110011" => q_unbuf <= my_rom(1203);
      when "0010010110100" => q_unbuf <= my_rom(1204);
      when "0010010110101" => q_unbuf <= my_rom(1205);
      when "0010010110110" => q_unbuf <= my_rom(1206);
      when "0010010110111" => q_unbuf <= my_rom(1207);
      when "0010010111000" => q_unbuf <= my_rom(1208);
      when "0010010111001" => q_unbuf <= my_rom(1209);
      when "0010010111010" => q_unbuf <= my_rom(1210);
      when "0010010111011" => q_unbuf <= my_rom(1211);
      when "0010010111100" => q_unbuf <= my_rom(1212);
      when "0010010111101" => q_unbuf <= my_rom(1213);
      when "0010010111110" => q_unbuf <= my_rom(1214);
      when "0010010111111" => q_unbuf <= my_rom(1215);
      when "0010011000000" => q_unbuf <= my_rom(1216);
      when "0010011000001" => q_unbuf <= my_rom(1217);
      when "0010011000010" => q_unbuf <= my_rom(1218);
      when "0010011000011" => q_unbuf <= my_rom(1219);
      when "0010011000100" => q_unbuf <= my_rom(1220);
      when "0010011000101" => q_unbuf <= my_rom(1221);
      when "0010011000110" => q_unbuf <= my_rom(1222);
      when "0010011000111" => q_unbuf <= my_rom(1223);
      when "0010011001000" => q_unbuf <= my_rom(1224);
      when "0010011001001" => q_unbuf <= my_rom(1225);
      when "0010011001010" => q_unbuf <= my_rom(1226);
      when "0010011001011" => q_unbuf <= my_rom(1227);
      when "0010011001100" => q_unbuf <= my_rom(1228);
      when "0010011001101" => q_unbuf <= my_rom(1229);
      when "0010011001110" => q_unbuf <= my_rom(1230);
      when "0010011001111" => q_unbuf <= my_rom(1231);
      when "0010011010000" => q_unbuf <= my_rom(1232);
      when "0010011010001" => q_unbuf <= my_rom(1233);
      when "0010011010010" => q_unbuf <= my_rom(1234);
      when "0010011010011" => q_unbuf <= my_rom(1235);
      when "0010011010100" => q_unbuf <= my_rom(1236);
      when "0010011010101" => q_unbuf <= my_rom(1237);
      when "0010011010110" => q_unbuf <= my_rom(1238);
      when "0010011010111" => q_unbuf <= my_rom(1239);
      when "0010011011000" => q_unbuf <= my_rom(1240);
      when "0010011011001" => q_unbuf <= my_rom(1241);
      when "0010011011010" => q_unbuf <= my_rom(1242);
      when "0010011011011" => q_unbuf <= my_rom(1243);
      when "0010011011100" => q_unbuf <= my_rom(1244);
      when "0010011011101" => q_unbuf <= my_rom(1245);
      when "0010011011110" => q_unbuf <= my_rom(1246);
      when "0010011011111" => q_unbuf <= my_rom(1247);
      when "0010011100000" => q_unbuf <= my_rom(1248);
      when "0010011100001" => q_unbuf <= my_rom(1249);
      when "0010011100010" => q_unbuf <= my_rom(1250);
      when "0010011100011" => q_unbuf <= my_rom(1251);
      when "0010011100100" => q_unbuf <= my_rom(1252);
      when "0010011100101" => q_unbuf <= my_rom(1253);
      when "0010011100110" => q_unbuf <= my_rom(1254);
      when "0010011100111" => q_unbuf <= my_rom(1255);
      when "0010011101000" => q_unbuf <= my_rom(1256);
      when "0010011101001" => q_unbuf <= my_rom(1257);
      when "0010011101010" => q_unbuf <= my_rom(1258);
      when "0010011101011" => q_unbuf <= my_rom(1259);
      when "0010011101100" => q_unbuf <= my_rom(1260);
      when "0010011101101" => q_unbuf <= my_rom(1261);
      when "0010011101110" => q_unbuf <= my_rom(1262);
      when "0010011101111" => q_unbuf <= my_rom(1263);
      when "0010011110000" => q_unbuf <= my_rom(1264);
      when "0010011110001" => q_unbuf <= my_rom(1265);
      when "0010011110010" => q_unbuf <= my_rom(1266);
      when "0010011110011" => q_unbuf <= my_rom(1267);
      when "0010011110100" => q_unbuf <= my_rom(1268);
      when "0010011110101" => q_unbuf <= my_rom(1269);
      when "0010011110110" => q_unbuf <= my_rom(1270);
      when "0010011110111" => q_unbuf <= my_rom(1271);
      when "0010011111000" => q_unbuf <= my_rom(1272);
      when "0010011111001" => q_unbuf <= my_rom(1273);
      when "0010011111010" => q_unbuf <= my_rom(1274);
      when "0010011111011" => q_unbuf <= my_rom(1275);
      when "0010011111100" => q_unbuf <= my_rom(1276);
      when "0010011111101" => q_unbuf <= my_rom(1277);
      when "0010011111110" => q_unbuf <= my_rom(1278);
      when "0010011111111" => q_unbuf <= my_rom(1279);
      when "0010100000000" => q_unbuf <= my_rom(1280);
      when "0010100000001" => q_unbuf <= my_rom(1281);
      when "0010100000010" => q_unbuf <= my_rom(1282);
      when "0010100000011" => q_unbuf <= my_rom(1283);
      when "0010100000100" => q_unbuf <= my_rom(1284);
      when "0010100000101" => q_unbuf <= my_rom(1285);
      when "0010100000110" => q_unbuf <= my_rom(1286);
      when "0010100000111" => q_unbuf <= my_rom(1287);
      when "0010100001000" => q_unbuf <= my_rom(1288);
      when "0010100001001" => q_unbuf <= my_rom(1289);
      when "0010100001010" => q_unbuf <= my_rom(1290);
      when "0010100001011" => q_unbuf <= my_rom(1291);
      when "0010100001100" => q_unbuf <= my_rom(1292);
      when "0010100001101" => q_unbuf <= my_rom(1293);
      when "0010100001110" => q_unbuf <= my_rom(1294);
      when "0010100001111" => q_unbuf <= my_rom(1295);
      when "0010100010000" => q_unbuf <= my_rom(1296);
      when "0010100010001" => q_unbuf <= my_rom(1297);
      when "0010100010010" => q_unbuf <= my_rom(1298);
      when "0010100010011" => q_unbuf <= my_rom(1299);
      when "0010100010100" => q_unbuf <= my_rom(1300);
      when "0010100010101" => q_unbuf <= my_rom(1301);
      when "0010100010110" => q_unbuf <= my_rom(1302);
      when "0010100010111" => q_unbuf <= my_rom(1303);
      when "0010100011000" => q_unbuf <= my_rom(1304);
      when "0010100011001" => q_unbuf <= my_rom(1305);
      when "0010100011010" => q_unbuf <= my_rom(1306);
      when "0010100011011" => q_unbuf <= my_rom(1307);
      when "0010100011100" => q_unbuf <= my_rom(1308);
      when "0010100011101" => q_unbuf <= my_rom(1309);
      when "0010100011110" => q_unbuf <= my_rom(1310);
      when "0010100011111" => q_unbuf <= my_rom(1311);
      when "0010100100000" => q_unbuf <= my_rom(1312);
      when "0010100100001" => q_unbuf <= my_rom(1313);
      when "0010100100010" => q_unbuf <= my_rom(1314);
      when "0010100100011" => q_unbuf <= my_rom(1315);
      when "0010100100100" => q_unbuf <= my_rom(1316);
      when "0010100100101" => q_unbuf <= my_rom(1317);
      when "0010100100110" => q_unbuf <= my_rom(1318);
      when "0010100100111" => q_unbuf <= my_rom(1319);
      when "0010100101000" => q_unbuf <= my_rom(1320);
      when "0010100101001" => q_unbuf <= my_rom(1321);
      when "0010100101010" => q_unbuf <= my_rom(1322);
      when "0010100101011" => q_unbuf <= my_rom(1323);
      when "0010100101100" => q_unbuf <= my_rom(1324);
      when "0010100101101" => q_unbuf <= my_rom(1325);
      when "0010100101110" => q_unbuf <= my_rom(1326);
      when "0010100101111" => q_unbuf <= my_rom(1327);
      when "0010100110000" => q_unbuf <= my_rom(1328);
      when "0010100110001" => q_unbuf <= my_rom(1329);
      when "0010100110010" => q_unbuf <= my_rom(1330);
      when "0010100110011" => q_unbuf <= my_rom(1331);
      when "0010100110100" => q_unbuf <= my_rom(1332);
      when "0010100110101" => q_unbuf <= my_rom(1333);
      when "0010100110110" => q_unbuf <= my_rom(1334);
      when "0010100110111" => q_unbuf <= my_rom(1335);
      when "0010100111000" => q_unbuf <= my_rom(1336);
      when "0010100111001" => q_unbuf <= my_rom(1337);
      when "0010100111010" => q_unbuf <= my_rom(1338);
      when "0010100111011" => q_unbuf <= my_rom(1339);
      when "0010100111100" => q_unbuf <= my_rom(1340);
      when "0010100111101" => q_unbuf <= my_rom(1341);
      when "0010100111110" => q_unbuf <= my_rom(1342);
      when "0010100111111" => q_unbuf <= my_rom(1343);
      when "0010101000000" => q_unbuf <= my_rom(1344);
      when "0010101000001" => q_unbuf <= my_rom(1345);
      when "0010101000010" => q_unbuf <= my_rom(1346);
      when "0010101000011" => q_unbuf <= my_rom(1347);
      when "0010101000100" => q_unbuf <= my_rom(1348);
      when "0010101000101" => q_unbuf <= my_rom(1349);
      when "0010101000110" => q_unbuf <= my_rom(1350);
      when "0010101000111" => q_unbuf <= my_rom(1351);
      when "0010101001000" => q_unbuf <= my_rom(1352);
      when "0010101001001" => q_unbuf <= my_rom(1353);
      when "0010101001010" => q_unbuf <= my_rom(1354);
      when "0010101001011" => q_unbuf <= my_rom(1355);
      when "0010101001100" => q_unbuf <= my_rom(1356);
      when "0010101001101" => q_unbuf <= my_rom(1357);
      when "0010101001110" => q_unbuf <= my_rom(1358);
      when "0010101001111" => q_unbuf <= my_rom(1359);
      when "0010101010000" => q_unbuf <= my_rom(1360);
      when "0010101010001" => q_unbuf <= my_rom(1361);
      when "0010101010010" => q_unbuf <= my_rom(1362);
      when "0010101010011" => q_unbuf <= my_rom(1363);
      when "0010101010100" => q_unbuf <= my_rom(1364);
      when "0010101010101" => q_unbuf <= my_rom(1365);
      when "0010101010110" => q_unbuf <= my_rom(1366);
      when "0010101010111" => q_unbuf <= my_rom(1367);
      when "0010101011000" => q_unbuf <= my_rom(1368);
      when "0010101011001" => q_unbuf <= my_rom(1369);
      when "0010101011010" => q_unbuf <= my_rom(1370);
      when "0010101011011" => q_unbuf <= my_rom(1371);
      when "0010101011100" => q_unbuf <= my_rom(1372);
      when "0010101011101" => q_unbuf <= my_rom(1373);
      when "0010101011110" => q_unbuf <= my_rom(1374);
      when "0010101011111" => q_unbuf <= my_rom(1375);
      when "0010101100000" => q_unbuf <= my_rom(1376);
      when "0010101100001" => q_unbuf <= my_rom(1377);
      when "0010101100010" => q_unbuf <= my_rom(1378);
      when "0010101100011" => q_unbuf <= my_rom(1379);
      when "0010101100100" => q_unbuf <= my_rom(1380);
      when "0010101100101" => q_unbuf <= my_rom(1381);
      when "0010101100110" => q_unbuf <= my_rom(1382);
      when "0010101100111" => q_unbuf <= my_rom(1383);
      when "0010101101000" => q_unbuf <= my_rom(1384);
      when "0010101101001" => q_unbuf <= my_rom(1385);
      when "0010101101010" => q_unbuf <= my_rom(1386);
      when "0010101101011" => q_unbuf <= my_rom(1387);
      when "0010101101100" => q_unbuf <= my_rom(1388);
      when "0010101101101" => q_unbuf <= my_rom(1389);
      when "0010101101110" => q_unbuf <= my_rom(1390);
      when "0010101101111" => q_unbuf <= my_rom(1391);
      when "0010101110000" => q_unbuf <= my_rom(1392);
      when "0010101110001" => q_unbuf <= my_rom(1393);
      when "0010101110010" => q_unbuf <= my_rom(1394);
      when "0010101110011" => q_unbuf <= my_rom(1395);
      when "0010101110100" => q_unbuf <= my_rom(1396);
      when "0010101110101" => q_unbuf <= my_rom(1397);
      when "0010101110110" => q_unbuf <= my_rom(1398);
      when "0010101110111" => q_unbuf <= my_rom(1399);
      when "0010101111000" => q_unbuf <= my_rom(1400);
      when "0010101111001" => q_unbuf <= my_rom(1401);
      when "0010101111010" => q_unbuf <= my_rom(1402);
      when "0010101111011" => q_unbuf <= my_rom(1403);
      when "0010101111100" => q_unbuf <= my_rom(1404);
      when "0010101111101" => q_unbuf <= my_rom(1405);
      when "0010101111110" => q_unbuf <= my_rom(1406);
      when "0010101111111" => q_unbuf <= my_rom(1407);
      when "0010110000000" => q_unbuf <= my_rom(1408);
      when "0010110000001" => q_unbuf <= my_rom(1409);
      when "0010110000010" => q_unbuf <= my_rom(1410);
      when "0010110000011" => q_unbuf <= my_rom(1411);
      when "0010110000100" => q_unbuf <= my_rom(1412);
      when "0010110000101" => q_unbuf <= my_rom(1413);
      when "0010110000110" => q_unbuf <= my_rom(1414);
      when "0010110000111" => q_unbuf <= my_rom(1415);
      when "0010110001000" => q_unbuf <= my_rom(1416);
      when "0010110001001" => q_unbuf <= my_rom(1417);
      when "0010110001010" => q_unbuf <= my_rom(1418);
      when "0010110001011" => q_unbuf <= my_rom(1419);
      when "0010110001100" => q_unbuf <= my_rom(1420);
      when "0010110001101" => q_unbuf <= my_rom(1421);
      when "0010110001110" => q_unbuf <= my_rom(1422);
      when "0010110001111" => q_unbuf <= my_rom(1423);
      when "0010110010000" => q_unbuf <= my_rom(1424);
      when "0010110010001" => q_unbuf <= my_rom(1425);
      when "0010110010010" => q_unbuf <= my_rom(1426);
      when "0010110010011" => q_unbuf <= my_rom(1427);
      when "0010110010100" => q_unbuf <= my_rom(1428);
      when "0010110010101" => q_unbuf <= my_rom(1429);
      when "0010110010110" => q_unbuf <= my_rom(1430);
      when "0010110010111" => q_unbuf <= my_rom(1431);
      when "0010110011000" => q_unbuf <= my_rom(1432);
      when "0010110011001" => q_unbuf <= my_rom(1433);
      when "0010110011010" => q_unbuf <= my_rom(1434);
      when "0010110011011" => q_unbuf <= my_rom(1435);
      when "0010110011100" => q_unbuf <= my_rom(1436);
      when "0010110011101" => q_unbuf <= my_rom(1437);
      when "0010110011110" => q_unbuf <= my_rom(1438);
      when "0010110011111" => q_unbuf <= my_rom(1439);
      when "0010110100000" => q_unbuf <= my_rom(1440);
      when "0010110100001" => q_unbuf <= my_rom(1441);
      when "0010110100010" => q_unbuf <= my_rom(1442);
      when "0010110100011" => q_unbuf <= my_rom(1443);
      when "0010110100100" => q_unbuf <= my_rom(1444);
      when "0010110100101" => q_unbuf <= my_rom(1445);
      when "0010110100110" => q_unbuf <= my_rom(1446);
      when "0010110100111" => q_unbuf <= my_rom(1447);
      when "0010110101000" => q_unbuf <= my_rom(1448);
      when "0010110101001" => q_unbuf <= my_rom(1449);
      when "0010110101010" => q_unbuf <= my_rom(1450);
      when "0010110101011" => q_unbuf <= my_rom(1451);
      when "0010110101100" => q_unbuf <= my_rom(1452);
      when "0010110101101" => q_unbuf <= my_rom(1453);
      when "0010110101110" => q_unbuf <= my_rom(1454);
      when "0010110101111" => q_unbuf <= my_rom(1455);
      when "0010110110000" => q_unbuf <= my_rom(1456);
      when "0010110110001" => q_unbuf <= my_rom(1457);
      when "0010110110010" => q_unbuf <= my_rom(1458);
      when "0010110110011" => q_unbuf <= my_rom(1459);
      when "0010110110100" => q_unbuf <= my_rom(1460);
      when "0010110110101" => q_unbuf <= my_rom(1461);
      when "0010110110110" => q_unbuf <= my_rom(1462);
      when "0010110110111" => q_unbuf <= my_rom(1463);
      when "0010110111000" => q_unbuf <= my_rom(1464);
      when "0010110111001" => q_unbuf <= my_rom(1465);
      when "0010110111010" => q_unbuf <= my_rom(1466);
      when "0010110111011" => q_unbuf <= my_rom(1467);
      when "0010110111100" => q_unbuf <= my_rom(1468);
      when "0010110111101" => q_unbuf <= my_rom(1469);
      when "0010110111110" => q_unbuf <= my_rom(1470);
      when "0010110111111" => q_unbuf <= my_rom(1471);
      when "0010111000000" => q_unbuf <= my_rom(1472);
      when "0010111000001" => q_unbuf <= my_rom(1473);
      when "0010111000010" => q_unbuf <= my_rom(1474);
      when "0010111000011" => q_unbuf <= my_rom(1475);
      when "0010111000100" => q_unbuf <= my_rom(1476);
      when "0010111000101" => q_unbuf <= my_rom(1477);
      when "0010111000110" => q_unbuf <= my_rom(1478);
      when "0010111000111" => q_unbuf <= my_rom(1479);
      when "0010111001000" => q_unbuf <= my_rom(1480);
      when "0010111001001" => q_unbuf <= my_rom(1481);
      when "0010111001010" => q_unbuf <= my_rom(1482);
      when "0010111001011" => q_unbuf <= my_rom(1483);
      when "0010111001100" => q_unbuf <= my_rom(1484);
      when "0010111001101" => q_unbuf <= my_rom(1485);
      when "0010111001110" => q_unbuf <= my_rom(1486);
      when "0010111001111" => q_unbuf <= my_rom(1487);
      when "0010111010000" => q_unbuf <= my_rom(1488);
      when "0010111010001" => q_unbuf <= my_rom(1489);
      when "0010111010010" => q_unbuf <= my_rom(1490);
      when "0010111010011" => q_unbuf <= my_rom(1491);
      when "0010111010100" => q_unbuf <= my_rom(1492);
      when "0010111010101" => q_unbuf <= my_rom(1493);
      when "0010111010110" => q_unbuf <= my_rom(1494);
      when "0010111010111" => q_unbuf <= my_rom(1495);
      when "0010111011000" => q_unbuf <= my_rom(1496);
      when "0010111011001" => q_unbuf <= my_rom(1497);
      when "0010111011010" => q_unbuf <= my_rom(1498);
      when "0010111011011" => q_unbuf <= my_rom(1499);
      when "0010111011100" => q_unbuf <= my_rom(1500);
      when "0010111011101" => q_unbuf <= my_rom(1501);
      when "0010111011110" => q_unbuf <= my_rom(1502);
      when "0010111011111" => q_unbuf <= my_rom(1503);
      when "0010111100000" => q_unbuf <= my_rom(1504);
      when "0010111100001" => q_unbuf <= my_rom(1505);
      when "0010111100010" => q_unbuf <= my_rom(1506);
      when "0010111100011" => q_unbuf <= my_rom(1507);
      when "0010111100100" => q_unbuf <= my_rom(1508);
      when "0010111100101" => q_unbuf <= my_rom(1509);
      when "0010111100110" => q_unbuf <= my_rom(1510);
      when "0010111100111" => q_unbuf <= my_rom(1511);
      when "0010111101000" => q_unbuf <= my_rom(1512);
      when "0010111101001" => q_unbuf <= my_rom(1513);
      when "0010111101010" => q_unbuf <= my_rom(1514);
      when "0010111101011" => q_unbuf <= my_rom(1515);
      when "0010111101100" => q_unbuf <= my_rom(1516);
      when "0010111101101" => q_unbuf <= my_rom(1517);
      when "0010111101110" => q_unbuf <= my_rom(1518);
      when "0010111101111" => q_unbuf <= my_rom(1519);
      when "0010111110000" => q_unbuf <= my_rom(1520);
      when "0010111110001" => q_unbuf <= my_rom(1521);
      when "0010111110010" => q_unbuf <= my_rom(1522);
      when "0010111110011" => q_unbuf <= my_rom(1523);
      when "0010111110100" => q_unbuf <= my_rom(1524);
      when "0010111110101" => q_unbuf <= my_rom(1525);
      when "0010111110110" => q_unbuf <= my_rom(1526);
      when "0010111110111" => q_unbuf <= my_rom(1527);
      when "0010111111000" => q_unbuf <= my_rom(1528);
      when "0010111111001" => q_unbuf <= my_rom(1529);
      when "0010111111010" => q_unbuf <= my_rom(1530);
      when "0010111111011" => q_unbuf <= my_rom(1531);
      when "0010111111100" => q_unbuf <= my_rom(1532);
      when "0010111111101" => q_unbuf <= my_rom(1533);
      when "0010111111110" => q_unbuf <= my_rom(1534);
      when "0010111111111" => q_unbuf <= my_rom(1535);
      when "0011000000000" => q_unbuf <= my_rom(1536);
      when "0011000000001" => q_unbuf <= my_rom(1537);
      when "0011000000010" => q_unbuf <= my_rom(1538);
      when "0011000000011" => q_unbuf <= my_rom(1539);
      when "0011000000100" => q_unbuf <= my_rom(1540);
      when "0011000000101" => q_unbuf <= my_rom(1541);
      when "0011000000110" => q_unbuf <= my_rom(1542);
      when "0011000000111" => q_unbuf <= my_rom(1543);
      when "0011000001000" => q_unbuf <= my_rom(1544);
      when "0011000001001" => q_unbuf <= my_rom(1545);
      when "0011000001010" => q_unbuf <= my_rom(1546);
      when "0011000001011" => q_unbuf <= my_rom(1547);
      when "0011000001100" => q_unbuf <= my_rom(1548);
      when "0011000001101" => q_unbuf <= my_rom(1549);
      when "0011000001110" => q_unbuf <= my_rom(1550);
      when "0011000001111" => q_unbuf <= my_rom(1551);
      when "0011000010000" => q_unbuf <= my_rom(1552);
      when "0011000010001" => q_unbuf <= my_rom(1553);
      when "0011000010010" => q_unbuf <= my_rom(1554);
      when "0011000010011" => q_unbuf <= my_rom(1555);
      when "0011000010100" => q_unbuf <= my_rom(1556);
      when "0011000010101" => q_unbuf <= my_rom(1557);
      when "0011000010110" => q_unbuf <= my_rom(1558);
      when "0011000010111" => q_unbuf <= my_rom(1559);
      when "0011000011000" => q_unbuf <= my_rom(1560);
      when "0011000011001" => q_unbuf <= my_rom(1561);
      when "0011000011010" => q_unbuf <= my_rom(1562);
      when "0011000011011" => q_unbuf <= my_rom(1563);
      when "0011000011100" => q_unbuf <= my_rom(1564);
      when "0011000011101" => q_unbuf <= my_rom(1565);
      when "0011000011110" => q_unbuf <= my_rom(1566);
      when "0011000011111" => q_unbuf <= my_rom(1567);
      when "0011000100000" => q_unbuf <= my_rom(1568);
      when "0011000100001" => q_unbuf <= my_rom(1569);
      when "0011000100010" => q_unbuf <= my_rom(1570);
      when "0011000100011" => q_unbuf <= my_rom(1571);
      when "0011000100100" => q_unbuf <= my_rom(1572);
      when "0011000100101" => q_unbuf <= my_rom(1573);
      when "0011000100110" => q_unbuf <= my_rom(1574);
      when "0011000100111" => q_unbuf <= my_rom(1575);
      when "0011000101000" => q_unbuf <= my_rom(1576);
      when "0011000101001" => q_unbuf <= my_rom(1577);
      when "0011000101010" => q_unbuf <= my_rom(1578);
      when "0011000101011" => q_unbuf <= my_rom(1579);
      when "0011000101100" => q_unbuf <= my_rom(1580);
      when "0011000101101" => q_unbuf <= my_rom(1581);
      when "0011000101110" => q_unbuf <= my_rom(1582);
      when "0011000101111" => q_unbuf <= my_rom(1583);
      when "0011000110000" => q_unbuf <= my_rom(1584);
      when "0011000110001" => q_unbuf <= my_rom(1585);
      when "0011000110010" => q_unbuf <= my_rom(1586);
      when "0011000110011" => q_unbuf <= my_rom(1587);
      when "0011000110100" => q_unbuf <= my_rom(1588);
      when "0011000110101" => q_unbuf <= my_rom(1589);
      when "0011000110110" => q_unbuf <= my_rom(1590);
      when "0011000110111" => q_unbuf <= my_rom(1591);
      when "0011000111000" => q_unbuf <= my_rom(1592);
      when "0011000111001" => q_unbuf <= my_rom(1593);
      when "0011000111010" => q_unbuf <= my_rom(1594);
      when "0011000111011" => q_unbuf <= my_rom(1595);
      when "0011000111100" => q_unbuf <= my_rom(1596);
      when "0011000111101" => q_unbuf <= my_rom(1597);
      when "0011000111110" => q_unbuf <= my_rom(1598);
      when "0011000111111" => q_unbuf <= my_rom(1599);
      when "0011001000000" => q_unbuf <= my_rom(1600);
      when "0011001000001" => q_unbuf <= my_rom(1601);
      when "0011001000010" => q_unbuf <= my_rom(1602);
      when "0011001000011" => q_unbuf <= my_rom(1603);
      when "0011001000100" => q_unbuf <= my_rom(1604);
      when "0011001000101" => q_unbuf <= my_rom(1605);
      when "0011001000110" => q_unbuf <= my_rom(1606);
      when "0011001000111" => q_unbuf <= my_rom(1607);
      when "0011001001000" => q_unbuf <= my_rom(1608);
      when "0011001001001" => q_unbuf <= my_rom(1609);
      when "0011001001010" => q_unbuf <= my_rom(1610);
      when "0011001001011" => q_unbuf <= my_rom(1611);
      when "0011001001100" => q_unbuf <= my_rom(1612);
      when "0011001001101" => q_unbuf <= my_rom(1613);
      when "0011001001110" => q_unbuf <= my_rom(1614);
      when "0011001001111" => q_unbuf <= my_rom(1615);
      when "0011001010000" => q_unbuf <= my_rom(1616);
      when "0011001010001" => q_unbuf <= my_rom(1617);
      when "0011001010010" => q_unbuf <= my_rom(1618);
      when "0011001010011" => q_unbuf <= my_rom(1619);
      when "0011001010100" => q_unbuf <= my_rom(1620);
      when "0011001010101" => q_unbuf <= my_rom(1621);
      when "0011001010110" => q_unbuf <= my_rom(1622);
      when "0011001010111" => q_unbuf <= my_rom(1623);
      when "0011001011000" => q_unbuf <= my_rom(1624);
      when "0011001011001" => q_unbuf <= my_rom(1625);
      when "0011001011010" => q_unbuf <= my_rom(1626);
      when "0011001011011" => q_unbuf <= my_rom(1627);
      when "0011001011100" => q_unbuf <= my_rom(1628);
      when "0011001011101" => q_unbuf <= my_rom(1629);
      when "0011001011110" => q_unbuf <= my_rom(1630);
      when "0011001011111" => q_unbuf <= my_rom(1631);
      when "0011001100000" => q_unbuf <= my_rom(1632);
      when "0011001100001" => q_unbuf <= my_rom(1633);
      when "0011001100010" => q_unbuf <= my_rom(1634);
      when "0011001100011" => q_unbuf <= my_rom(1635);
      when "0011001100100" => q_unbuf <= my_rom(1636);
      when "0011001100101" => q_unbuf <= my_rom(1637);
      when "0011001100110" => q_unbuf <= my_rom(1638);
      when "0011001100111" => q_unbuf <= my_rom(1639);
      when "0011001101000" => q_unbuf <= my_rom(1640);
      when "0011001101001" => q_unbuf <= my_rom(1641);
      when "0011001101010" => q_unbuf <= my_rom(1642);
      when "0011001101011" => q_unbuf <= my_rom(1643);
      when "0011001101100" => q_unbuf <= my_rom(1644);
      when "0011001101101" => q_unbuf <= my_rom(1645);
      when "0011001101110" => q_unbuf <= my_rom(1646);
      when "0011001101111" => q_unbuf <= my_rom(1647);
      when "0011001110000" => q_unbuf <= my_rom(1648);
      when "0011001110001" => q_unbuf <= my_rom(1649);
      when "0011001110010" => q_unbuf <= my_rom(1650);
      when "0011001110011" => q_unbuf <= my_rom(1651);
      when "0011001110100" => q_unbuf <= my_rom(1652);
      when "0011001110101" => q_unbuf <= my_rom(1653);
      when "0011001110110" => q_unbuf <= my_rom(1654);
      when "0011001110111" => q_unbuf <= my_rom(1655);
      when "0011001111000" => q_unbuf <= my_rom(1656);
      when "0011001111001" => q_unbuf <= my_rom(1657);
      when "0011001111010" => q_unbuf <= my_rom(1658);
      when "0011001111011" => q_unbuf <= my_rom(1659);
      when "0011001111100" => q_unbuf <= my_rom(1660);
      when "0011001111101" => q_unbuf <= my_rom(1661);
      when "0011001111110" => q_unbuf <= my_rom(1662);
      when "0011001111111" => q_unbuf <= my_rom(1663);
      when "0011010000000" => q_unbuf <= my_rom(1664);
      when "0011010000001" => q_unbuf <= my_rom(1665);
      when "0011010000010" => q_unbuf <= my_rom(1666);
      when "0011010000011" => q_unbuf <= my_rom(1667);
      when "0011010000100" => q_unbuf <= my_rom(1668);
      when "0011010000101" => q_unbuf <= my_rom(1669);
      when "0011010000110" => q_unbuf <= my_rom(1670);
      when "0011010000111" => q_unbuf <= my_rom(1671);
      when "0011010001000" => q_unbuf <= my_rom(1672);
      when "0011010001001" => q_unbuf <= my_rom(1673);
      when "0011010001010" => q_unbuf <= my_rom(1674);
      when "0011010001011" => q_unbuf <= my_rom(1675);
      when "0011010001100" => q_unbuf <= my_rom(1676);
      when "0011010001101" => q_unbuf <= my_rom(1677);
      when "0011010001110" => q_unbuf <= my_rom(1678);
      when "0011010001111" => q_unbuf <= my_rom(1679);
      when "0011010010000" => q_unbuf <= my_rom(1680);
      when "0011010010001" => q_unbuf <= my_rom(1681);
      when "0011010010010" => q_unbuf <= my_rom(1682);
      when "0011010010011" => q_unbuf <= my_rom(1683);
      when "0011010010100" => q_unbuf <= my_rom(1684);
      when "0011010010101" => q_unbuf <= my_rom(1685);
      when "0011010010110" => q_unbuf <= my_rom(1686);
      when "0011010010111" => q_unbuf <= my_rom(1687);
      when "0011010011000" => q_unbuf <= my_rom(1688);
      when "0011010011001" => q_unbuf <= my_rom(1689);
      when "0011010011010" => q_unbuf <= my_rom(1690);
      when "0011010011011" => q_unbuf <= my_rom(1691);
      when "0011010011100" => q_unbuf <= my_rom(1692);
      when "0011010011101" => q_unbuf <= my_rom(1693);
      when "0011010011110" => q_unbuf <= my_rom(1694);
      when "0011010011111" => q_unbuf <= my_rom(1695);
      when "0011010100000" => q_unbuf <= my_rom(1696);
      when "0011010100001" => q_unbuf <= my_rom(1697);
      when "0011010100010" => q_unbuf <= my_rom(1698);
      when "0011010100011" => q_unbuf <= my_rom(1699);
      when "0011010100100" => q_unbuf <= my_rom(1700);
      when "0011010100101" => q_unbuf <= my_rom(1701);
      when "0011010100110" => q_unbuf <= my_rom(1702);
      when "0011010100111" => q_unbuf <= my_rom(1703);
      when "0011010101000" => q_unbuf <= my_rom(1704);
      when "0011010101001" => q_unbuf <= my_rom(1705);
      when "0011010101010" => q_unbuf <= my_rom(1706);
      when "0011010101011" => q_unbuf <= my_rom(1707);
      when "0011010101100" => q_unbuf <= my_rom(1708);
      when "0011010101101" => q_unbuf <= my_rom(1709);
      when "0011010101110" => q_unbuf <= my_rom(1710);
      when "0011010101111" => q_unbuf <= my_rom(1711);
      when "0011010110000" => q_unbuf <= my_rom(1712);
      when "0011010110001" => q_unbuf <= my_rom(1713);
      when "0011010110010" => q_unbuf <= my_rom(1714);
      when "0011010110011" => q_unbuf <= my_rom(1715);
      when "0011010110100" => q_unbuf <= my_rom(1716);
      when "0011010110101" => q_unbuf <= my_rom(1717);
      when "0011010110110" => q_unbuf <= my_rom(1718);
      when "0011010110111" => q_unbuf <= my_rom(1719);
      when "0011010111000" => q_unbuf <= my_rom(1720);
      when "0011010111001" => q_unbuf <= my_rom(1721);
      when "0011010111010" => q_unbuf <= my_rom(1722);
      when "0011010111011" => q_unbuf <= my_rom(1723);
      when "0011010111100" => q_unbuf <= my_rom(1724);
      when "0011010111101" => q_unbuf <= my_rom(1725);
      when "0011010111110" => q_unbuf <= my_rom(1726);
      when "0011010111111" => q_unbuf <= my_rom(1727);
      when "0011011000000" => q_unbuf <= my_rom(1728);
      when "0011011000001" => q_unbuf <= my_rom(1729);
      when "0011011000010" => q_unbuf <= my_rom(1730);
      when "0011011000011" => q_unbuf <= my_rom(1731);
      when "0011011000100" => q_unbuf <= my_rom(1732);
      when "0011011000101" => q_unbuf <= my_rom(1733);
      when "0011011000110" => q_unbuf <= my_rom(1734);
      when "0011011000111" => q_unbuf <= my_rom(1735);
      when "0011011001000" => q_unbuf <= my_rom(1736);
      when "0011011001001" => q_unbuf <= my_rom(1737);
      when "0011011001010" => q_unbuf <= my_rom(1738);
      when "0011011001011" => q_unbuf <= my_rom(1739);
      when "0011011001100" => q_unbuf <= my_rom(1740);
      when "0011011001101" => q_unbuf <= my_rom(1741);
      when "0011011001110" => q_unbuf <= my_rom(1742);
      when "0011011001111" => q_unbuf <= my_rom(1743);
      when "0011011010000" => q_unbuf <= my_rom(1744);
      when "0011011010001" => q_unbuf <= my_rom(1745);
      when "0011011010010" => q_unbuf <= my_rom(1746);
      when "0011011010011" => q_unbuf <= my_rom(1747);
      when "0011011010100" => q_unbuf <= my_rom(1748);
      when "0011011010101" => q_unbuf <= my_rom(1749);
      when "0011011010110" => q_unbuf <= my_rom(1750);
      when "0011011010111" => q_unbuf <= my_rom(1751);
      when "0011011011000" => q_unbuf <= my_rom(1752);
      when "0011011011001" => q_unbuf <= my_rom(1753);
      when "0011011011010" => q_unbuf <= my_rom(1754);
      when "0011011011011" => q_unbuf <= my_rom(1755);
      when "0011011011100" => q_unbuf <= my_rom(1756);
      when "0011011011101" => q_unbuf <= my_rom(1757);
      when "0011011011110" => q_unbuf <= my_rom(1758);
      when "0011011011111" => q_unbuf <= my_rom(1759);
      when "0011011100000" => q_unbuf <= my_rom(1760);
      when "0011011100001" => q_unbuf <= my_rom(1761);
      when "0011011100010" => q_unbuf <= my_rom(1762);
      when "0011011100011" => q_unbuf <= my_rom(1763);
      when "0011011100100" => q_unbuf <= my_rom(1764);
      when "0011011100101" => q_unbuf <= my_rom(1765);
      when "0011011100110" => q_unbuf <= my_rom(1766);
      when "0011011100111" => q_unbuf <= my_rom(1767);
      when "0011011101000" => q_unbuf <= my_rom(1768);
      when "0011011101001" => q_unbuf <= my_rom(1769);
      when "0011011101010" => q_unbuf <= my_rom(1770);
      when "0011011101011" => q_unbuf <= my_rom(1771);
      when "0011011101100" => q_unbuf <= my_rom(1772);
      when "0011011101101" => q_unbuf <= my_rom(1773);
      when "0011011101110" => q_unbuf <= my_rom(1774);
      when "0011011101111" => q_unbuf <= my_rom(1775);
      when "0011011110000" => q_unbuf <= my_rom(1776);
      when "0011011110001" => q_unbuf <= my_rom(1777);
      when "0011011110010" => q_unbuf <= my_rom(1778);
      when "0011011110011" => q_unbuf <= my_rom(1779);
      when "0011011110100" => q_unbuf <= my_rom(1780);
      when "0011011110101" => q_unbuf <= my_rom(1781);
      when "0011011110110" => q_unbuf <= my_rom(1782);
      when "0011011110111" => q_unbuf <= my_rom(1783);
      when "0011011111000" => q_unbuf <= my_rom(1784);
      when "0011011111001" => q_unbuf <= my_rom(1785);
      when "0011011111010" => q_unbuf <= my_rom(1786);
      when "0011011111011" => q_unbuf <= my_rom(1787);
      when "0011011111100" => q_unbuf <= my_rom(1788);
      when "0011011111101" => q_unbuf <= my_rom(1789);
      when "0011011111110" => q_unbuf <= my_rom(1790);
      when "0011011111111" => q_unbuf <= my_rom(1791);
      when "0011100000000" => q_unbuf <= my_rom(1792);
      when "0011100000001" => q_unbuf <= my_rom(1793);
      when "0011100000010" => q_unbuf <= my_rom(1794);
      when "0011100000011" => q_unbuf <= my_rom(1795);
      when "0011100000100" => q_unbuf <= my_rom(1796);
      when "0011100000101" => q_unbuf <= my_rom(1797);
      when "0011100000110" => q_unbuf <= my_rom(1798);
      when "0011100000111" => q_unbuf <= my_rom(1799);
      when "0011100001000" => q_unbuf <= my_rom(1800);
      when "0011100001001" => q_unbuf <= my_rom(1801);
      when "0011100001010" => q_unbuf <= my_rom(1802);
      when "0011100001011" => q_unbuf <= my_rom(1803);
      when "0011100001100" => q_unbuf <= my_rom(1804);
      when "0011100001101" => q_unbuf <= my_rom(1805);
      when "0011100001110" => q_unbuf <= my_rom(1806);
      when "0011100001111" => q_unbuf <= my_rom(1807);
      when "0011100010000" => q_unbuf <= my_rom(1808);
      when "0011100010001" => q_unbuf <= my_rom(1809);
      when "0011100010010" => q_unbuf <= my_rom(1810);
      when "0011100010011" => q_unbuf <= my_rom(1811);
      when "0011100010100" => q_unbuf <= my_rom(1812);
      when "0011100010101" => q_unbuf <= my_rom(1813);
      when "0011100010110" => q_unbuf <= my_rom(1814);
      when "0011100010111" => q_unbuf <= my_rom(1815);
      when "0011100011000" => q_unbuf <= my_rom(1816);
      when "0011100011001" => q_unbuf <= my_rom(1817);
      when "0011100011010" => q_unbuf <= my_rom(1818);
      when "0011100011011" => q_unbuf <= my_rom(1819);
      when "0011100011100" => q_unbuf <= my_rom(1820);
      when "0011100011101" => q_unbuf <= my_rom(1821);
      when "0011100011110" => q_unbuf <= my_rom(1822);
      when "0011100011111" => q_unbuf <= my_rom(1823);
      when "0011100100000" => q_unbuf <= my_rom(1824);
      when "0011100100001" => q_unbuf <= my_rom(1825);
      when "0011100100010" => q_unbuf <= my_rom(1826);
      when "0011100100011" => q_unbuf <= my_rom(1827);
      when "0011100100100" => q_unbuf <= my_rom(1828);
      when "0011100100101" => q_unbuf <= my_rom(1829);
      when "0011100100110" => q_unbuf <= my_rom(1830);
      when "0011100100111" => q_unbuf <= my_rom(1831);
      when "0011100101000" => q_unbuf <= my_rom(1832);
      when "0011100101001" => q_unbuf <= my_rom(1833);
      when "0011100101010" => q_unbuf <= my_rom(1834);
      when "0011100101011" => q_unbuf <= my_rom(1835);
      when "0011100101100" => q_unbuf <= my_rom(1836);
      when "0011100101101" => q_unbuf <= my_rom(1837);
      when "0011100101110" => q_unbuf <= my_rom(1838);
      when "0011100101111" => q_unbuf <= my_rom(1839);
      when "0011100110000" => q_unbuf <= my_rom(1840);
      when "0011100110001" => q_unbuf <= my_rom(1841);
      when "0011100110010" => q_unbuf <= my_rom(1842);
      when "0011100110011" => q_unbuf <= my_rom(1843);
      when "0011100110100" => q_unbuf <= my_rom(1844);
      when "0011100110101" => q_unbuf <= my_rom(1845);
      when "0011100110110" => q_unbuf <= my_rom(1846);
      when "0011100110111" => q_unbuf <= my_rom(1847);
      when "0011100111000" => q_unbuf <= my_rom(1848);
      when "0011100111001" => q_unbuf <= my_rom(1849);
      when "0011100111010" => q_unbuf <= my_rom(1850);
      when "0011100111011" => q_unbuf <= my_rom(1851);
      when "0011100111100" => q_unbuf <= my_rom(1852);
      when "0011100111101" => q_unbuf <= my_rom(1853);
      when "0011100111110" => q_unbuf <= my_rom(1854);
      when "0011100111111" => q_unbuf <= my_rom(1855);
      when "0011101000000" => q_unbuf <= my_rom(1856);
      when "0011101000001" => q_unbuf <= my_rom(1857);
      when "0011101000010" => q_unbuf <= my_rom(1858);
      when "0011101000011" => q_unbuf <= my_rom(1859);
      when "0011101000100" => q_unbuf <= my_rom(1860);
      when "0011101000101" => q_unbuf <= my_rom(1861);
      when "0011101000110" => q_unbuf <= my_rom(1862);
      when "0011101000111" => q_unbuf <= my_rom(1863);
      when "0011101001000" => q_unbuf <= my_rom(1864);
      when "0011101001001" => q_unbuf <= my_rom(1865);
      when "0011101001010" => q_unbuf <= my_rom(1866);
      when "0011101001011" => q_unbuf <= my_rom(1867);
      when "0011101001100" => q_unbuf <= my_rom(1868);
      when "0011101001101" => q_unbuf <= my_rom(1869);
      when "0011101001110" => q_unbuf <= my_rom(1870);
      when "0011101001111" => q_unbuf <= my_rom(1871);
      when "0011101010000" => q_unbuf <= my_rom(1872);
      when "0011101010001" => q_unbuf <= my_rom(1873);
      when "0011101010010" => q_unbuf <= my_rom(1874);
      when "0011101010011" => q_unbuf <= my_rom(1875);
      when "0011101010100" => q_unbuf <= my_rom(1876);
      when "0011101010101" => q_unbuf <= my_rom(1877);
      when "0011101010110" => q_unbuf <= my_rom(1878);
      when "0011101010111" => q_unbuf <= my_rom(1879);
      when "0011101011000" => q_unbuf <= my_rom(1880);
      when "0011101011001" => q_unbuf <= my_rom(1881);
      when "0011101011010" => q_unbuf <= my_rom(1882);
      when "0011101011011" => q_unbuf <= my_rom(1883);
      when "0011101011100" => q_unbuf <= my_rom(1884);
      when "0011101011101" => q_unbuf <= my_rom(1885);
      when "0011101011110" => q_unbuf <= my_rom(1886);
      when "0011101011111" => q_unbuf <= my_rom(1887);
      when "0011101100000" => q_unbuf <= my_rom(1888);
      when "0011101100001" => q_unbuf <= my_rom(1889);
      when "0011101100010" => q_unbuf <= my_rom(1890);
      when "0011101100011" => q_unbuf <= my_rom(1891);
      when "0011101100100" => q_unbuf <= my_rom(1892);
      when "0011101100101" => q_unbuf <= my_rom(1893);
      when "0011101100110" => q_unbuf <= my_rom(1894);
      when "0011101100111" => q_unbuf <= my_rom(1895);
      when "0011101101000" => q_unbuf <= my_rom(1896);
      when "0011101101001" => q_unbuf <= my_rom(1897);
      when "0011101101010" => q_unbuf <= my_rom(1898);
      when "0011101101011" => q_unbuf <= my_rom(1899);
      when "0011101101100" => q_unbuf <= my_rom(1900);
      when "0011101101101" => q_unbuf <= my_rom(1901);
      when "0011101101110" => q_unbuf <= my_rom(1902);
      when "0011101101111" => q_unbuf <= my_rom(1903);
      when "0011101110000" => q_unbuf <= my_rom(1904);
      when "0011101110001" => q_unbuf <= my_rom(1905);
      when "0011101110010" => q_unbuf <= my_rom(1906);
      when "0011101110011" => q_unbuf <= my_rom(1907);
      when "0011101110100" => q_unbuf <= my_rom(1908);
      when "0011101110101" => q_unbuf <= my_rom(1909);
      when "0011101110110" => q_unbuf <= my_rom(1910);
      when "0011101110111" => q_unbuf <= my_rom(1911);
      when "0011101111000" => q_unbuf <= my_rom(1912);
      when "0011101111001" => q_unbuf <= my_rom(1913);
      when "0011101111010" => q_unbuf <= my_rom(1914);
      when "0011101111011" => q_unbuf <= my_rom(1915);
      when "0011101111100" => q_unbuf <= my_rom(1916);
      when "0011101111101" => q_unbuf <= my_rom(1917);
      when "0011101111110" => q_unbuf <= my_rom(1918);
      when "0011101111111" => q_unbuf <= my_rom(1919);
      when "0011110000000" => q_unbuf <= my_rom(1920);
      when "0011110000001" => q_unbuf <= my_rom(1921);
      when "0011110000010" => q_unbuf <= my_rom(1922);
      when "0011110000011" => q_unbuf <= my_rom(1923);
      when "0011110000100" => q_unbuf <= my_rom(1924);
      when "0011110000101" => q_unbuf <= my_rom(1925);
      when "0011110000110" => q_unbuf <= my_rom(1926);
      when "0011110000111" => q_unbuf <= my_rom(1927);
      when "0011110001000" => q_unbuf <= my_rom(1928);
      when "0011110001001" => q_unbuf <= my_rom(1929);
      when "0011110001010" => q_unbuf <= my_rom(1930);
      when "0011110001011" => q_unbuf <= my_rom(1931);
      when "0011110001100" => q_unbuf <= my_rom(1932);
      when "0011110001101" => q_unbuf <= my_rom(1933);
      when "0011110001110" => q_unbuf <= my_rom(1934);
      when "0011110001111" => q_unbuf <= my_rom(1935);
      when "0011110010000" => q_unbuf <= my_rom(1936);
      when "0011110010001" => q_unbuf <= my_rom(1937);
      when "0011110010010" => q_unbuf <= my_rom(1938);
      when "0011110010011" => q_unbuf <= my_rom(1939);
      when "0011110010100" => q_unbuf <= my_rom(1940);
      when "0011110010101" => q_unbuf <= my_rom(1941);
      when "0011110010110" => q_unbuf <= my_rom(1942);
      when "0011110010111" => q_unbuf <= my_rom(1943);
      when "0011110011000" => q_unbuf <= my_rom(1944);
      when "0011110011001" => q_unbuf <= my_rom(1945);
      when "0011110011010" => q_unbuf <= my_rom(1946);
      when "0011110011011" => q_unbuf <= my_rom(1947);
      when "0011110011100" => q_unbuf <= my_rom(1948);
      when "0011110011101" => q_unbuf <= my_rom(1949);
      when "0011110011110" => q_unbuf <= my_rom(1950);
      when "0011110011111" => q_unbuf <= my_rom(1951);
      when "0011110100000" => q_unbuf <= my_rom(1952);
      when "0011110100001" => q_unbuf <= my_rom(1953);
      when "0011110100010" => q_unbuf <= my_rom(1954);
      when "0011110100011" => q_unbuf <= my_rom(1955);
      when "0011110100100" => q_unbuf <= my_rom(1956);
      when "0011110100101" => q_unbuf <= my_rom(1957);
      when "0011110100110" => q_unbuf <= my_rom(1958);
      when "0011110100111" => q_unbuf <= my_rom(1959);
      when "0011110101000" => q_unbuf <= my_rom(1960);
      when "0011110101001" => q_unbuf <= my_rom(1961);
      when "0011110101010" => q_unbuf <= my_rom(1962);
      when "0011110101011" => q_unbuf <= my_rom(1963);
      when "0011110101100" => q_unbuf <= my_rom(1964);
      when "0011110101101" => q_unbuf <= my_rom(1965);
      when "0011110101110" => q_unbuf <= my_rom(1966);
      when "0011110101111" => q_unbuf <= my_rom(1967);
      when "0011110110000" => q_unbuf <= my_rom(1968);
      when "0011110110001" => q_unbuf <= my_rom(1969);
      when "0011110110010" => q_unbuf <= my_rom(1970);
      when "0011110110011" => q_unbuf <= my_rom(1971);
      when "0011110110100" => q_unbuf <= my_rom(1972);
      when "0011110110101" => q_unbuf <= my_rom(1973);
      when "0011110110110" => q_unbuf <= my_rom(1974);
      when "0011110110111" => q_unbuf <= my_rom(1975);
      when "0011110111000" => q_unbuf <= my_rom(1976);
      when "0011110111001" => q_unbuf <= my_rom(1977);
      when "0011110111010" => q_unbuf <= my_rom(1978);
      when "0011110111011" => q_unbuf <= my_rom(1979);
      when "0011110111100" => q_unbuf <= my_rom(1980);
      when "0011110111101" => q_unbuf <= my_rom(1981);
      when "0011110111110" => q_unbuf <= my_rom(1982);
      when "0011110111111" => q_unbuf <= my_rom(1983);
      when "0011111000000" => q_unbuf <= my_rom(1984);
      when "0011111000001" => q_unbuf <= my_rom(1985);
      when "0011111000010" => q_unbuf <= my_rom(1986);
      when "0011111000011" => q_unbuf <= my_rom(1987);
      when "0011111000100" => q_unbuf <= my_rom(1988);
      when "0011111000101" => q_unbuf <= my_rom(1989);
      when "0011111000110" => q_unbuf <= my_rom(1990);
      when "0011111000111" => q_unbuf <= my_rom(1991);
      when "0011111001000" => q_unbuf <= my_rom(1992);
      when "0011111001001" => q_unbuf <= my_rom(1993);
      when "0011111001010" => q_unbuf <= my_rom(1994);
      when "0011111001011" => q_unbuf <= my_rom(1995);
      when "0011111001100" => q_unbuf <= my_rom(1996);
      when "0011111001101" => q_unbuf <= my_rom(1997);
      when "0011111001110" => q_unbuf <= my_rom(1998);
      when "0011111001111" => q_unbuf <= my_rom(1999);
      when "0011111010000" => q_unbuf <= my_rom(2000);
      when "0011111010001" => q_unbuf <= my_rom(2001);
      when "0011111010010" => q_unbuf <= my_rom(2002);
      when "0011111010011" => q_unbuf <= my_rom(2003);
      when "0011111010100" => q_unbuf <= my_rom(2004);
      when "0011111010101" => q_unbuf <= my_rom(2005);
      when "0011111010110" => q_unbuf <= my_rom(2006);
      when "0011111010111" => q_unbuf <= my_rom(2007);
      when "0011111011000" => q_unbuf <= my_rom(2008);
      when "0011111011001" => q_unbuf <= my_rom(2009);
      when "0011111011010" => q_unbuf <= my_rom(2010);
      when "0011111011011" => q_unbuf <= my_rom(2011);
      when "0011111011100" => q_unbuf <= my_rom(2012);
      when "0011111011101" => q_unbuf <= my_rom(2013);
      when "0011111011110" => q_unbuf <= my_rom(2014);
      when "0011111011111" => q_unbuf <= my_rom(2015);
      when "0011111100000" => q_unbuf <= my_rom(2016);
      when "0011111100001" => q_unbuf <= my_rom(2017);
      when "0011111100010" => q_unbuf <= my_rom(2018);
      when "0011111100011" => q_unbuf <= my_rom(2019);
      when "0011111100100" => q_unbuf <= my_rom(2020);
      when "0011111100101" => q_unbuf <= my_rom(2021);
      when "0011111100110" => q_unbuf <= my_rom(2022);
      when "0011111100111" => q_unbuf <= my_rom(2023);
      when "0011111101000" => q_unbuf <= my_rom(2024);
      when "0011111101001" => q_unbuf <= my_rom(2025);
      when "0011111101010" => q_unbuf <= my_rom(2026);
      when "0011111101011" => q_unbuf <= my_rom(2027);
      when "0011111101100" => q_unbuf <= my_rom(2028);
      when "0011111101101" => q_unbuf <= my_rom(2029);
      when "0011111101110" => q_unbuf <= my_rom(2030);
      when "0011111101111" => q_unbuf <= my_rom(2031);
      when "0011111110000" => q_unbuf <= my_rom(2032);
      when "0011111110001" => q_unbuf <= my_rom(2033);
      when "0011111110010" => q_unbuf <= my_rom(2034);
      when "0011111110011" => q_unbuf <= my_rom(2035);
      when "0011111110100" => q_unbuf <= my_rom(2036);
      when "0011111110101" => q_unbuf <= my_rom(2037);
      when "0011111110110" => q_unbuf <= my_rom(2038);
      when "0011111110111" => q_unbuf <= my_rom(2039);
      when "0011111111000" => q_unbuf <= my_rom(2040);
      when "0011111111001" => q_unbuf <= my_rom(2041);
      when "0011111111010" => q_unbuf <= my_rom(2042);
      when "0011111111011" => q_unbuf <= my_rom(2043);
      when "0011111111100" => q_unbuf <= my_rom(2044);
      when "0011111111101" => q_unbuf <= my_rom(2045);
      when "0011111111110" => q_unbuf <= my_rom(2046);
      when "0011111111111" => q_unbuf <= my_rom(2047);
      when "0100000000000" => q_unbuf <= my_rom(2048);
      when "0100000000001" => q_unbuf <= my_rom(2049);
      when "0100000000010" => q_unbuf <= my_rom(2050);
      when "0100000000011" => q_unbuf <= my_rom(2051);
      when "0100000000100" => q_unbuf <= my_rom(2052);
      when "0100000000101" => q_unbuf <= my_rom(2053);
      when "0100000000110" => q_unbuf <= my_rom(2054);
      when "0100000000111" => q_unbuf <= my_rom(2055);
      when "0100000001000" => q_unbuf <= my_rom(2056);
      when "0100000001001" => q_unbuf <= my_rom(2057);
      when "0100000001010" => q_unbuf <= my_rom(2058);
      when "0100000001011" => q_unbuf <= my_rom(2059);
      when "0100000001100" => q_unbuf <= my_rom(2060);
      when "0100000001101" => q_unbuf <= my_rom(2061);
      when "0100000001110" => q_unbuf <= my_rom(2062);
      when "0100000001111" => q_unbuf <= my_rom(2063);
      when "0100000010000" => q_unbuf <= my_rom(2064);
      when "0100000010001" => q_unbuf <= my_rom(2065);
      when "0100000010010" => q_unbuf <= my_rom(2066);
      when "0100000010011" => q_unbuf <= my_rom(2067);
      when "0100000010100" => q_unbuf <= my_rom(2068);
      when "0100000010101" => q_unbuf <= my_rom(2069);
      when "0100000010110" => q_unbuf <= my_rom(2070);
      when "0100000010111" => q_unbuf <= my_rom(2071);
      when "0100000011000" => q_unbuf <= my_rom(2072);
      when "0100000011001" => q_unbuf <= my_rom(2073);
      when "0100000011010" => q_unbuf <= my_rom(2074);
      when "0100000011011" => q_unbuf <= my_rom(2075);
      when "0100000011100" => q_unbuf <= my_rom(2076);
      when "0100000011101" => q_unbuf <= my_rom(2077);
      when "0100000011110" => q_unbuf <= my_rom(2078);
      when "0100000011111" => q_unbuf <= my_rom(2079);
      when "0100000100000" => q_unbuf <= my_rom(2080);
      when "0100000100001" => q_unbuf <= my_rom(2081);
      when "0100000100010" => q_unbuf <= my_rom(2082);
      when "0100000100011" => q_unbuf <= my_rom(2083);
      when "0100000100100" => q_unbuf <= my_rom(2084);
      when "0100000100101" => q_unbuf <= my_rom(2085);
      when "0100000100110" => q_unbuf <= my_rom(2086);
      when "0100000100111" => q_unbuf <= my_rom(2087);
      when "0100000101000" => q_unbuf <= my_rom(2088);
      when "0100000101001" => q_unbuf <= my_rom(2089);
      when "0100000101010" => q_unbuf <= my_rom(2090);
      when "0100000101011" => q_unbuf <= my_rom(2091);
      when "0100000101100" => q_unbuf <= my_rom(2092);
      when "0100000101101" => q_unbuf <= my_rom(2093);
      when "0100000101110" => q_unbuf <= my_rom(2094);
      when "0100000101111" => q_unbuf <= my_rom(2095);
      when "0100000110000" => q_unbuf <= my_rom(2096);
      when "0100000110001" => q_unbuf <= my_rom(2097);
      when "0100000110010" => q_unbuf <= my_rom(2098);
      when "0100000110011" => q_unbuf <= my_rom(2099);
      when "0100000110100" => q_unbuf <= my_rom(2100);
      when "0100000110101" => q_unbuf <= my_rom(2101);
      when "0100000110110" => q_unbuf <= my_rom(2102);
      when "0100000110111" => q_unbuf <= my_rom(2103);
      when "0100000111000" => q_unbuf <= my_rom(2104);
      when "0100000111001" => q_unbuf <= my_rom(2105);
      when "0100000111010" => q_unbuf <= my_rom(2106);
      when "0100000111011" => q_unbuf <= my_rom(2107);
      when "0100000111100" => q_unbuf <= my_rom(2108);
      when "0100000111101" => q_unbuf <= my_rom(2109);
      when "0100000111110" => q_unbuf <= my_rom(2110);
      when "0100000111111" => q_unbuf <= my_rom(2111);
      when "0100001000000" => q_unbuf <= my_rom(2112);
      when "0100001000001" => q_unbuf <= my_rom(2113);
      when "0100001000010" => q_unbuf <= my_rom(2114);
      when "0100001000011" => q_unbuf <= my_rom(2115);
      when "0100001000100" => q_unbuf <= my_rom(2116);
      when "0100001000101" => q_unbuf <= my_rom(2117);
      when "0100001000110" => q_unbuf <= my_rom(2118);
      when "0100001000111" => q_unbuf <= my_rom(2119);
      when "0100001001000" => q_unbuf <= my_rom(2120);
      when "0100001001001" => q_unbuf <= my_rom(2121);
      when "0100001001010" => q_unbuf <= my_rom(2122);
      when "0100001001011" => q_unbuf <= my_rom(2123);
      when "0100001001100" => q_unbuf <= my_rom(2124);
      when "0100001001101" => q_unbuf <= my_rom(2125);
      when "0100001001110" => q_unbuf <= my_rom(2126);
      when "0100001001111" => q_unbuf <= my_rom(2127);
      when "0100001010000" => q_unbuf <= my_rom(2128);
      when "0100001010001" => q_unbuf <= my_rom(2129);
      when "0100001010010" => q_unbuf <= my_rom(2130);
      when "0100001010011" => q_unbuf <= my_rom(2131);
      when "0100001010100" => q_unbuf <= my_rom(2132);
      when "0100001010101" => q_unbuf <= my_rom(2133);
      when "0100001010110" => q_unbuf <= my_rom(2134);
      when "0100001010111" => q_unbuf <= my_rom(2135);
      when "0100001011000" => q_unbuf <= my_rom(2136);
      when "0100001011001" => q_unbuf <= my_rom(2137);
      when "0100001011010" => q_unbuf <= my_rom(2138);
      when "0100001011011" => q_unbuf <= my_rom(2139);
      when "0100001011100" => q_unbuf <= my_rom(2140);
      when "0100001011101" => q_unbuf <= my_rom(2141);
      when "0100001011110" => q_unbuf <= my_rom(2142);
      when "0100001011111" => q_unbuf <= my_rom(2143);
      when "0100001100000" => q_unbuf <= my_rom(2144);
      when "0100001100001" => q_unbuf <= my_rom(2145);
      when "0100001100010" => q_unbuf <= my_rom(2146);
      when "0100001100011" => q_unbuf <= my_rom(2147);
      when "0100001100100" => q_unbuf <= my_rom(2148);
      when "0100001100101" => q_unbuf <= my_rom(2149);
      when "0100001100110" => q_unbuf <= my_rom(2150);
      when "0100001100111" => q_unbuf <= my_rom(2151);
      when "0100001101000" => q_unbuf <= my_rom(2152);
      when "0100001101001" => q_unbuf <= my_rom(2153);
      when "0100001101010" => q_unbuf <= my_rom(2154);
      when "0100001101011" => q_unbuf <= my_rom(2155);
      when "0100001101100" => q_unbuf <= my_rom(2156);
      when "0100001101101" => q_unbuf <= my_rom(2157);
      when "0100001101110" => q_unbuf <= my_rom(2158);
      when "0100001101111" => q_unbuf <= my_rom(2159);
      when "0100001110000" => q_unbuf <= my_rom(2160);
      when "0100001110001" => q_unbuf <= my_rom(2161);
      when "0100001110010" => q_unbuf <= my_rom(2162);
      when "0100001110011" => q_unbuf <= my_rom(2163);
      when "0100001110100" => q_unbuf <= my_rom(2164);
      when "0100001110101" => q_unbuf <= my_rom(2165);
      when "0100001110110" => q_unbuf <= my_rom(2166);
      when "0100001110111" => q_unbuf <= my_rom(2167);
      when "0100001111000" => q_unbuf <= my_rom(2168);
      when "0100001111001" => q_unbuf <= my_rom(2169);
      when "0100001111010" => q_unbuf <= my_rom(2170);
      when "0100001111011" => q_unbuf <= my_rom(2171);
      when "0100001111100" => q_unbuf <= my_rom(2172);
      when "0100001111101" => q_unbuf <= my_rom(2173);
      when "0100001111110" => q_unbuf <= my_rom(2174);
      when "0100001111111" => q_unbuf <= my_rom(2175);
      when "0100010000000" => q_unbuf <= my_rom(2176);
      when "0100010000001" => q_unbuf <= my_rom(2177);
      when "0100010000010" => q_unbuf <= my_rom(2178);
      when "0100010000011" => q_unbuf <= my_rom(2179);
      when "0100010000100" => q_unbuf <= my_rom(2180);
      when "0100010000101" => q_unbuf <= my_rom(2181);
      when "0100010000110" => q_unbuf <= my_rom(2182);
      when "0100010000111" => q_unbuf <= my_rom(2183);
      when "0100010001000" => q_unbuf <= my_rom(2184);
      when "0100010001001" => q_unbuf <= my_rom(2185);
      when "0100010001010" => q_unbuf <= my_rom(2186);
      when "0100010001011" => q_unbuf <= my_rom(2187);
      when "0100010001100" => q_unbuf <= my_rom(2188);
      when "0100010001101" => q_unbuf <= my_rom(2189);
      when "0100010001110" => q_unbuf <= my_rom(2190);
      when "0100010001111" => q_unbuf <= my_rom(2191);
      when "0100010010000" => q_unbuf <= my_rom(2192);
      when "0100010010001" => q_unbuf <= my_rom(2193);
      when "0100010010010" => q_unbuf <= my_rom(2194);
      when "0100010010011" => q_unbuf <= my_rom(2195);
      when "0100010010100" => q_unbuf <= my_rom(2196);
      when "0100010010101" => q_unbuf <= my_rom(2197);
      when "0100010010110" => q_unbuf <= my_rom(2198);
      when "0100010010111" => q_unbuf <= my_rom(2199);
      when "0100010011000" => q_unbuf <= my_rom(2200);
      when "0100010011001" => q_unbuf <= my_rom(2201);
      when "0100010011010" => q_unbuf <= my_rom(2202);
      when "0100010011011" => q_unbuf <= my_rom(2203);
      when "0100010011100" => q_unbuf <= my_rom(2204);
      when "0100010011101" => q_unbuf <= my_rom(2205);
      when "0100010011110" => q_unbuf <= my_rom(2206);
      when "0100010011111" => q_unbuf <= my_rom(2207);
      when "0100010100000" => q_unbuf <= my_rom(2208);
      when "0100010100001" => q_unbuf <= my_rom(2209);
      when "0100010100010" => q_unbuf <= my_rom(2210);
      when "0100010100011" => q_unbuf <= my_rom(2211);
      when "0100010100100" => q_unbuf <= my_rom(2212);
      when "0100010100101" => q_unbuf <= my_rom(2213);
      when "0100010100110" => q_unbuf <= my_rom(2214);
      when "0100010100111" => q_unbuf <= my_rom(2215);
      when "0100010101000" => q_unbuf <= my_rom(2216);
      when "0100010101001" => q_unbuf <= my_rom(2217);
      when "0100010101010" => q_unbuf <= my_rom(2218);
      when "0100010101011" => q_unbuf <= my_rom(2219);
      when "0100010101100" => q_unbuf <= my_rom(2220);
      when "0100010101101" => q_unbuf <= my_rom(2221);
      when "0100010101110" => q_unbuf <= my_rom(2222);
      when "0100010101111" => q_unbuf <= my_rom(2223);
      when "0100010110000" => q_unbuf <= my_rom(2224);
      when "0100010110001" => q_unbuf <= my_rom(2225);
      when "0100010110010" => q_unbuf <= my_rom(2226);
      when "0100010110011" => q_unbuf <= my_rom(2227);
      when "0100010110100" => q_unbuf <= my_rom(2228);
      when "0100010110101" => q_unbuf <= my_rom(2229);
      when "0100010110110" => q_unbuf <= my_rom(2230);
      when "0100010110111" => q_unbuf <= my_rom(2231);
      when "0100010111000" => q_unbuf <= my_rom(2232);
      when "0100010111001" => q_unbuf <= my_rom(2233);
      when "0100010111010" => q_unbuf <= my_rom(2234);
      when "0100010111011" => q_unbuf <= my_rom(2235);
      when "0100010111100" => q_unbuf <= my_rom(2236);
      when "0100010111101" => q_unbuf <= my_rom(2237);
      when "0100010111110" => q_unbuf <= my_rom(2238);
      when "0100010111111" => q_unbuf <= my_rom(2239);
      when "0100011000000" => q_unbuf <= my_rom(2240);
      when "0100011000001" => q_unbuf <= my_rom(2241);
      when "0100011000010" => q_unbuf <= my_rom(2242);
      when "0100011000011" => q_unbuf <= my_rom(2243);
      when "0100011000100" => q_unbuf <= my_rom(2244);
      when "0100011000101" => q_unbuf <= my_rom(2245);
      when "0100011000110" => q_unbuf <= my_rom(2246);
      when "0100011000111" => q_unbuf <= my_rom(2247);
      when "0100011001000" => q_unbuf <= my_rom(2248);
      when "0100011001001" => q_unbuf <= my_rom(2249);
      when "0100011001010" => q_unbuf <= my_rom(2250);
      when "0100011001011" => q_unbuf <= my_rom(2251);
      when "0100011001100" => q_unbuf <= my_rom(2252);
      when "0100011001101" => q_unbuf <= my_rom(2253);
      when "0100011001110" => q_unbuf <= my_rom(2254);
      when "0100011001111" => q_unbuf <= my_rom(2255);
      when "0100011010000" => q_unbuf <= my_rom(2256);
      when "0100011010001" => q_unbuf <= my_rom(2257);
      when "0100011010010" => q_unbuf <= my_rom(2258);
      when "0100011010011" => q_unbuf <= my_rom(2259);
      when "0100011010100" => q_unbuf <= my_rom(2260);
      when "0100011010101" => q_unbuf <= my_rom(2261);
      when "0100011010110" => q_unbuf <= my_rom(2262);
      when "0100011010111" => q_unbuf <= my_rom(2263);
      when "0100011011000" => q_unbuf <= my_rom(2264);
      when "0100011011001" => q_unbuf <= my_rom(2265);
      when "0100011011010" => q_unbuf <= my_rom(2266);
      when "0100011011011" => q_unbuf <= my_rom(2267);
      when "0100011011100" => q_unbuf <= my_rom(2268);
      when "0100011011101" => q_unbuf <= my_rom(2269);
      when "0100011011110" => q_unbuf <= my_rom(2270);
      when "0100011011111" => q_unbuf <= my_rom(2271);
      when "0100011100000" => q_unbuf <= my_rom(2272);
      when "0100011100001" => q_unbuf <= my_rom(2273);
      when "0100011100010" => q_unbuf <= my_rom(2274);
      when "0100011100011" => q_unbuf <= my_rom(2275);
      when "0100011100100" => q_unbuf <= my_rom(2276);
      when "0100011100101" => q_unbuf <= my_rom(2277);
      when "0100011100110" => q_unbuf <= my_rom(2278);
      when "0100011100111" => q_unbuf <= my_rom(2279);
      when "0100011101000" => q_unbuf <= my_rom(2280);
      when "0100011101001" => q_unbuf <= my_rom(2281);
      when "0100011101010" => q_unbuf <= my_rom(2282);
      when "0100011101011" => q_unbuf <= my_rom(2283);
      when "0100011101100" => q_unbuf <= my_rom(2284);
      when "0100011101101" => q_unbuf <= my_rom(2285);
      when "0100011101110" => q_unbuf <= my_rom(2286);
      when "0100011101111" => q_unbuf <= my_rom(2287);
      when "0100011110000" => q_unbuf <= my_rom(2288);
      when "0100011110001" => q_unbuf <= my_rom(2289);
      when "0100011110010" => q_unbuf <= my_rom(2290);
      when "0100011110011" => q_unbuf <= my_rom(2291);
      when "0100011110100" => q_unbuf <= my_rom(2292);
      when "0100011110101" => q_unbuf <= my_rom(2293);
      when "0100011110110" => q_unbuf <= my_rom(2294);
      when "0100011110111" => q_unbuf <= my_rom(2295);
      when "0100011111000" => q_unbuf <= my_rom(2296);
      when "0100011111001" => q_unbuf <= my_rom(2297);
      when "0100011111010" => q_unbuf <= my_rom(2298);
      when "0100011111011" => q_unbuf <= my_rom(2299);
      when "0100011111100" => q_unbuf <= my_rom(2300);
      when "0100011111101" => q_unbuf <= my_rom(2301);
      when "0100011111110" => q_unbuf <= my_rom(2302);
      when "0100011111111" => q_unbuf <= my_rom(2303);
      when "0100100000000" => q_unbuf <= my_rom(2304);
      when "0100100000001" => q_unbuf <= my_rom(2305);
      when "0100100000010" => q_unbuf <= my_rom(2306);
      when "0100100000011" => q_unbuf <= my_rom(2307);
      when "0100100000100" => q_unbuf <= my_rom(2308);
      when "0100100000101" => q_unbuf <= my_rom(2309);
      when "0100100000110" => q_unbuf <= my_rom(2310);
      when "0100100000111" => q_unbuf <= my_rom(2311);
      when "0100100001000" => q_unbuf <= my_rom(2312);
      when "0100100001001" => q_unbuf <= my_rom(2313);
      when "0100100001010" => q_unbuf <= my_rom(2314);
      when "0100100001011" => q_unbuf <= my_rom(2315);
      when "0100100001100" => q_unbuf <= my_rom(2316);
      when "0100100001101" => q_unbuf <= my_rom(2317);
      when "0100100001110" => q_unbuf <= my_rom(2318);
      when "0100100001111" => q_unbuf <= my_rom(2319);
      when "0100100010000" => q_unbuf <= my_rom(2320);
      when "0100100010001" => q_unbuf <= my_rom(2321);
      when "0100100010010" => q_unbuf <= my_rom(2322);
      when "0100100010011" => q_unbuf <= my_rom(2323);
      when "0100100010100" => q_unbuf <= my_rom(2324);
      when "0100100010101" => q_unbuf <= my_rom(2325);
      when "0100100010110" => q_unbuf <= my_rom(2326);
      when "0100100010111" => q_unbuf <= my_rom(2327);
      when "0100100011000" => q_unbuf <= my_rom(2328);
      when "0100100011001" => q_unbuf <= my_rom(2329);
      when "0100100011010" => q_unbuf <= my_rom(2330);
      when "0100100011011" => q_unbuf <= my_rom(2331);
      when "0100100011100" => q_unbuf <= my_rom(2332);
      when "0100100011101" => q_unbuf <= my_rom(2333);
      when "0100100011110" => q_unbuf <= my_rom(2334);
      when "0100100011111" => q_unbuf <= my_rom(2335);
      when "0100100100000" => q_unbuf <= my_rom(2336);
      when "0100100100001" => q_unbuf <= my_rom(2337);
      when "0100100100010" => q_unbuf <= my_rom(2338);
      when "0100100100011" => q_unbuf <= my_rom(2339);
      when "0100100100100" => q_unbuf <= my_rom(2340);
      when "0100100100101" => q_unbuf <= my_rom(2341);
      when "0100100100110" => q_unbuf <= my_rom(2342);
      when "0100100100111" => q_unbuf <= my_rom(2343);
      when "0100100101000" => q_unbuf <= my_rom(2344);
      when "0100100101001" => q_unbuf <= my_rom(2345);
      when "0100100101010" => q_unbuf <= my_rom(2346);
      when "0100100101011" => q_unbuf <= my_rom(2347);
      when "0100100101100" => q_unbuf <= my_rom(2348);
      when "0100100101101" => q_unbuf <= my_rom(2349);
      when "0100100101110" => q_unbuf <= my_rom(2350);
      when "0100100101111" => q_unbuf <= my_rom(2351);
      when "0100100110000" => q_unbuf <= my_rom(2352);
      when "0100100110001" => q_unbuf <= my_rom(2353);
      when "0100100110010" => q_unbuf <= my_rom(2354);
      when "0100100110011" => q_unbuf <= my_rom(2355);
      when "0100100110100" => q_unbuf <= my_rom(2356);
      when "0100100110101" => q_unbuf <= my_rom(2357);
      when "0100100110110" => q_unbuf <= my_rom(2358);
      when "0100100110111" => q_unbuf <= my_rom(2359);
      when "0100100111000" => q_unbuf <= my_rom(2360);
      when "0100100111001" => q_unbuf <= my_rom(2361);
      when "0100100111010" => q_unbuf <= my_rom(2362);
      when "0100100111011" => q_unbuf <= my_rom(2363);
      when "0100100111100" => q_unbuf <= my_rom(2364);
      when "0100100111101" => q_unbuf <= my_rom(2365);
      when "0100100111110" => q_unbuf <= my_rom(2366);
      when "0100100111111" => q_unbuf <= my_rom(2367);
      when "0100101000000" => q_unbuf <= my_rom(2368);
      when "0100101000001" => q_unbuf <= my_rom(2369);
      when "0100101000010" => q_unbuf <= my_rom(2370);
      when "0100101000011" => q_unbuf <= my_rom(2371);
      when "0100101000100" => q_unbuf <= my_rom(2372);
      when "0100101000101" => q_unbuf <= my_rom(2373);
      when "0100101000110" => q_unbuf <= my_rom(2374);
      when "0100101000111" => q_unbuf <= my_rom(2375);
      when "0100101001000" => q_unbuf <= my_rom(2376);
      when "0100101001001" => q_unbuf <= my_rom(2377);
      when "0100101001010" => q_unbuf <= my_rom(2378);
      when "0100101001011" => q_unbuf <= my_rom(2379);
      when "0100101001100" => q_unbuf <= my_rom(2380);
      when "0100101001101" => q_unbuf <= my_rom(2381);
      when "0100101001110" => q_unbuf <= my_rom(2382);
      when "0100101001111" => q_unbuf <= my_rom(2383);
      when "0100101010000" => q_unbuf <= my_rom(2384);
      when "0100101010001" => q_unbuf <= my_rom(2385);
      when "0100101010010" => q_unbuf <= my_rom(2386);
      when "0100101010011" => q_unbuf <= my_rom(2387);
      when "0100101010100" => q_unbuf <= my_rom(2388);
      when "0100101010101" => q_unbuf <= my_rom(2389);
      when "0100101010110" => q_unbuf <= my_rom(2390);
      when "0100101010111" => q_unbuf <= my_rom(2391);
      when "0100101011000" => q_unbuf <= my_rom(2392);
      when "0100101011001" => q_unbuf <= my_rom(2393);
      when "0100101011010" => q_unbuf <= my_rom(2394);
      when "0100101011011" => q_unbuf <= my_rom(2395);
      when "0100101011100" => q_unbuf <= my_rom(2396);
      when "0100101011101" => q_unbuf <= my_rom(2397);
      when "0100101011110" => q_unbuf <= my_rom(2398);
      when "0100101011111" => q_unbuf <= my_rom(2399);
      when "0100101100000" => q_unbuf <= my_rom(2400);
      when "0100101100001" => q_unbuf <= my_rom(2401);
      when "0100101100010" => q_unbuf <= my_rom(2402);
      when "0100101100011" => q_unbuf <= my_rom(2403);
      when "0100101100100" => q_unbuf <= my_rom(2404);
      when "0100101100101" => q_unbuf <= my_rom(2405);
      when "0100101100110" => q_unbuf <= my_rom(2406);
      when "0100101100111" => q_unbuf <= my_rom(2407);
      when "0100101101000" => q_unbuf <= my_rom(2408);
      when "0100101101001" => q_unbuf <= my_rom(2409);
      when "0100101101010" => q_unbuf <= my_rom(2410);
      when "0100101101011" => q_unbuf <= my_rom(2411);
      when "0100101101100" => q_unbuf <= my_rom(2412);
      when "0100101101101" => q_unbuf <= my_rom(2413);
      when "0100101101110" => q_unbuf <= my_rom(2414);
      when "0100101101111" => q_unbuf <= my_rom(2415);
      when "0100101110000" => q_unbuf <= my_rom(2416);
      when "0100101110001" => q_unbuf <= my_rom(2417);
      when "0100101110010" => q_unbuf <= my_rom(2418);
      when "0100101110011" => q_unbuf <= my_rom(2419);
      when "0100101110100" => q_unbuf <= my_rom(2420);
      when "0100101110101" => q_unbuf <= my_rom(2421);
      when "0100101110110" => q_unbuf <= my_rom(2422);
      when "0100101110111" => q_unbuf <= my_rom(2423);
      when "0100101111000" => q_unbuf <= my_rom(2424);
      when "0100101111001" => q_unbuf <= my_rom(2425);
      when "0100101111010" => q_unbuf <= my_rom(2426);
      when "0100101111011" => q_unbuf <= my_rom(2427);
      when "0100101111100" => q_unbuf <= my_rom(2428);
      when "0100101111101" => q_unbuf <= my_rom(2429);
      when "0100101111110" => q_unbuf <= my_rom(2430);
      when "0100101111111" => q_unbuf <= my_rom(2431);
      when "0100110000000" => q_unbuf <= my_rom(2432);
      when "0100110000001" => q_unbuf <= my_rom(2433);
      when "0100110000010" => q_unbuf <= my_rom(2434);
      when "0100110000011" => q_unbuf <= my_rom(2435);
      when "0100110000100" => q_unbuf <= my_rom(2436);
      when "0100110000101" => q_unbuf <= my_rom(2437);
      when "0100110000110" => q_unbuf <= my_rom(2438);
      when "0100110000111" => q_unbuf <= my_rom(2439);
      when "0100110001000" => q_unbuf <= my_rom(2440);
      when "0100110001001" => q_unbuf <= my_rom(2441);
      when "0100110001010" => q_unbuf <= my_rom(2442);
      when "0100110001011" => q_unbuf <= my_rom(2443);
      when "0100110001100" => q_unbuf <= my_rom(2444);
      when "0100110001101" => q_unbuf <= my_rom(2445);
      when "0100110001110" => q_unbuf <= my_rom(2446);
      when "0100110001111" => q_unbuf <= my_rom(2447);
      when "0100110010000" => q_unbuf <= my_rom(2448);
      when "0100110010001" => q_unbuf <= my_rom(2449);
      when "0100110010010" => q_unbuf <= my_rom(2450);
      when "0100110010011" => q_unbuf <= my_rom(2451);
      when "0100110010100" => q_unbuf <= my_rom(2452);
      when "0100110010101" => q_unbuf <= my_rom(2453);
      when "0100110010110" => q_unbuf <= my_rom(2454);
      when "0100110010111" => q_unbuf <= my_rom(2455);
      when "0100110011000" => q_unbuf <= my_rom(2456);
      when "0100110011001" => q_unbuf <= my_rom(2457);
      when "0100110011010" => q_unbuf <= my_rom(2458);
      when "0100110011011" => q_unbuf <= my_rom(2459);
      when "0100110011100" => q_unbuf <= my_rom(2460);
      when "0100110011101" => q_unbuf <= my_rom(2461);
      when "0100110011110" => q_unbuf <= my_rom(2462);
      when "0100110011111" => q_unbuf <= my_rom(2463);
      when "0100110100000" => q_unbuf <= my_rom(2464);
      when "0100110100001" => q_unbuf <= my_rom(2465);
      when "0100110100010" => q_unbuf <= my_rom(2466);
      when "0100110100011" => q_unbuf <= my_rom(2467);
      when "0100110100100" => q_unbuf <= my_rom(2468);
      when "0100110100101" => q_unbuf <= my_rom(2469);
      when "0100110100110" => q_unbuf <= my_rom(2470);
      when "0100110100111" => q_unbuf <= my_rom(2471);
      when "0100110101000" => q_unbuf <= my_rom(2472);
      when "0100110101001" => q_unbuf <= my_rom(2473);
      when "0100110101010" => q_unbuf <= my_rom(2474);
      when "0100110101011" => q_unbuf <= my_rom(2475);
      when "0100110101100" => q_unbuf <= my_rom(2476);
      when "0100110101101" => q_unbuf <= my_rom(2477);
      when "0100110101110" => q_unbuf <= my_rom(2478);
      when "0100110101111" => q_unbuf <= my_rom(2479);
      when "0100110110000" => q_unbuf <= my_rom(2480);
      when "0100110110001" => q_unbuf <= my_rom(2481);
      when "0100110110010" => q_unbuf <= my_rom(2482);
      when "0100110110011" => q_unbuf <= my_rom(2483);
      when "0100110110100" => q_unbuf <= my_rom(2484);
      when "0100110110101" => q_unbuf <= my_rom(2485);
      when "0100110110110" => q_unbuf <= my_rom(2486);
      when "0100110110111" => q_unbuf <= my_rom(2487);
      when "0100110111000" => q_unbuf <= my_rom(2488);
      when "0100110111001" => q_unbuf <= my_rom(2489);
      when "0100110111010" => q_unbuf <= my_rom(2490);
      when "0100110111011" => q_unbuf <= my_rom(2491);
      when "0100110111100" => q_unbuf <= my_rom(2492);
      when "0100110111101" => q_unbuf <= my_rom(2493);
      when "0100110111110" => q_unbuf <= my_rom(2494);
      when "0100110111111" => q_unbuf <= my_rom(2495);
      when "0100111000000" => q_unbuf <= my_rom(2496);
      when "0100111000001" => q_unbuf <= my_rom(2497);
      when "0100111000010" => q_unbuf <= my_rom(2498);
      when "0100111000011" => q_unbuf <= my_rom(2499);
      when "0100111000100" => q_unbuf <= my_rom(2500);
      when "0100111000101" => q_unbuf <= my_rom(2501);
      when "0100111000110" => q_unbuf <= my_rom(2502);
      when "0100111000111" => q_unbuf <= my_rom(2503);
      when "0100111001000" => q_unbuf <= my_rom(2504);
      when "0100111001001" => q_unbuf <= my_rom(2505);
      when "0100111001010" => q_unbuf <= my_rom(2506);
      when "0100111001011" => q_unbuf <= my_rom(2507);
      when "0100111001100" => q_unbuf <= my_rom(2508);
      when "0100111001101" => q_unbuf <= my_rom(2509);
      when "0100111001110" => q_unbuf <= my_rom(2510);
      when "0100111001111" => q_unbuf <= my_rom(2511);
      when "0100111010000" => q_unbuf <= my_rom(2512);
      when "0100111010001" => q_unbuf <= my_rom(2513);
      when "0100111010010" => q_unbuf <= my_rom(2514);
      when "0100111010011" => q_unbuf <= my_rom(2515);
      when "0100111010100" => q_unbuf <= my_rom(2516);
      when "0100111010101" => q_unbuf <= my_rom(2517);
      when "0100111010110" => q_unbuf <= my_rom(2518);
      when "0100111010111" => q_unbuf <= my_rom(2519);
      when "0100111011000" => q_unbuf <= my_rom(2520);
      when "0100111011001" => q_unbuf <= my_rom(2521);
      when "0100111011010" => q_unbuf <= my_rom(2522);
      when "0100111011011" => q_unbuf <= my_rom(2523);
      when "0100111011100" => q_unbuf <= my_rom(2524);
      when "0100111011101" => q_unbuf <= my_rom(2525);
      when "0100111011110" => q_unbuf <= my_rom(2526);
      when "0100111011111" => q_unbuf <= my_rom(2527);
      when "0100111100000" => q_unbuf <= my_rom(2528);
      when "0100111100001" => q_unbuf <= my_rom(2529);
      when "0100111100010" => q_unbuf <= my_rom(2530);
      when "0100111100011" => q_unbuf <= my_rom(2531);
      when "0100111100100" => q_unbuf <= my_rom(2532);
      when "0100111100101" => q_unbuf <= my_rom(2533);
      when "0100111100110" => q_unbuf <= my_rom(2534);
      when "0100111100111" => q_unbuf <= my_rom(2535);
      when "0100111101000" => q_unbuf <= my_rom(2536);
      when "0100111101001" => q_unbuf <= my_rom(2537);
      when "0100111101010" => q_unbuf <= my_rom(2538);
      when "0100111101011" => q_unbuf <= my_rom(2539);
      when "0100111101100" => q_unbuf <= my_rom(2540);
      when "0100111101101" => q_unbuf <= my_rom(2541);
      when "0100111101110" => q_unbuf <= my_rom(2542);
      when "0100111101111" => q_unbuf <= my_rom(2543);
      when "0100111110000" => q_unbuf <= my_rom(2544);
      when "0100111110001" => q_unbuf <= my_rom(2545);
      when "0100111110010" => q_unbuf <= my_rom(2546);
      when "0100111110011" => q_unbuf <= my_rom(2547);
      when "0100111110100" => q_unbuf <= my_rom(2548);
      when "0100111110101" => q_unbuf <= my_rom(2549);
      when "0100111110110" => q_unbuf <= my_rom(2550);
      when "0100111110111" => q_unbuf <= my_rom(2551);
      when "0100111111000" => q_unbuf <= my_rom(2552);
      when "0100111111001" => q_unbuf <= my_rom(2553);
      when "0100111111010" => q_unbuf <= my_rom(2554);
      when "0100111111011" => q_unbuf <= my_rom(2555);
      when "0100111111100" => q_unbuf <= my_rom(2556);
      when "0100111111101" => q_unbuf <= my_rom(2557);
      when "0100111111110" => q_unbuf <= my_rom(2558);
      when "0100111111111" => q_unbuf <= my_rom(2559);
      when "0101000000000" => q_unbuf <= my_rom(2560);
      when "0101000000001" => q_unbuf <= my_rom(2561);
      when "0101000000010" => q_unbuf <= my_rom(2562);
      when "0101000000011" => q_unbuf <= my_rom(2563);
      when "0101000000100" => q_unbuf <= my_rom(2564);
      when "0101000000101" => q_unbuf <= my_rom(2565);
      when "0101000000110" => q_unbuf <= my_rom(2566);
      when "0101000000111" => q_unbuf <= my_rom(2567);
      when "0101000001000" => q_unbuf <= my_rom(2568);
      when "0101000001001" => q_unbuf <= my_rom(2569);
      when "0101000001010" => q_unbuf <= my_rom(2570);
      when "0101000001011" => q_unbuf <= my_rom(2571);
      when "0101000001100" => q_unbuf <= my_rom(2572);
      when "0101000001101" => q_unbuf <= my_rom(2573);
      when "0101000001110" => q_unbuf <= my_rom(2574);
      when "0101000001111" => q_unbuf <= my_rom(2575);
      when "0101000010000" => q_unbuf <= my_rom(2576);
      when "0101000010001" => q_unbuf <= my_rom(2577);
      when "0101000010010" => q_unbuf <= my_rom(2578);
      when "0101000010011" => q_unbuf <= my_rom(2579);
      when "0101000010100" => q_unbuf <= my_rom(2580);
      when "0101000010101" => q_unbuf <= my_rom(2581);
      when "0101000010110" => q_unbuf <= my_rom(2582);
      when "0101000010111" => q_unbuf <= my_rom(2583);
      when "0101000011000" => q_unbuf <= my_rom(2584);
      when "0101000011001" => q_unbuf <= my_rom(2585);
      when "0101000011010" => q_unbuf <= my_rom(2586);
      when "0101000011011" => q_unbuf <= my_rom(2587);
      when "0101000011100" => q_unbuf <= my_rom(2588);
      when "0101000011101" => q_unbuf <= my_rom(2589);
      when "0101000011110" => q_unbuf <= my_rom(2590);
      when "0101000011111" => q_unbuf <= my_rom(2591);
      when "0101000100000" => q_unbuf <= my_rom(2592);
      when "0101000100001" => q_unbuf <= my_rom(2593);
      when "0101000100010" => q_unbuf <= my_rom(2594);
      when "0101000100011" => q_unbuf <= my_rom(2595);
      when "0101000100100" => q_unbuf <= my_rom(2596);
      when "0101000100101" => q_unbuf <= my_rom(2597);
      when "0101000100110" => q_unbuf <= my_rom(2598);
      when "0101000100111" => q_unbuf <= my_rom(2599);
      when "0101000101000" => q_unbuf <= my_rom(2600);
      when "0101000101001" => q_unbuf <= my_rom(2601);
      when "0101000101010" => q_unbuf <= my_rom(2602);
      when "0101000101011" => q_unbuf <= my_rom(2603);
      when "0101000101100" => q_unbuf <= my_rom(2604);
      when "0101000101101" => q_unbuf <= my_rom(2605);
      when "0101000101110" => q_unbuf <= my_rom(2606);
      when "0101000101111" => q_unbuf <= my_rom(2607);
      when "0101000110000" => q_unbuf <= my_rom(2608);
      when "0101000110001" => q_unbuf <= my_rom(2609);
      when "0101000110010" => q_unbuf <= my_rom(2610);
      when "0101000110011" => q_unbuf <= my_rom(2611);
      when "0101000110100" => q_unbuf <= my_rom(2612);
      when "0101000110101" => q_unbuf <= my_rom(2613);
      when "0101000110110" => q_unbuf <= my_rom(2614);
      when "0101000110111" => q_unbuf <= my_rom(2615);
      when "0101000111000" => q_unbuf <= my_rom(2616);
      when "0101000111001" => q_unbuf <= my_rom(2617);
      when "0101000111010" => q_unbuf <= my_rom(2618);
      when "0101000111011" => q_unbuf <= my_rom(2619);
      when "0101000111100" => q_unbuf <= my_rom(2620);
      when "0101000111101" => q_unbuf <= my_rom(2621);
      when "0101000111110" => q_unbuf <= my_rom(2622);
      when "0101000111111" => q_unbuf <= my_rom(2623);
      when "0101001000000" => q_unbuf <= my_rom(2624);
      when "0101001000001" => q_unbuf <= my_rom(2625);
      when "0101001000010" => q_unbuf <= my_rom(2626);
      when "0101001000011" => q_unbuf <= my_rom(2627);
      when "0101001000100" => q_unbuf <= my_rom(2628);
      when "0101001000101" => q_unbuf <= my_rom(2629);
      when "0101001000110" => q_unbuf <= my_rom(2630);
      when "0101001000111" => q_unbuf <= my_rom(2631);
      when "0101001001000" => q_unbuf <= my_rom(2632);
      when "0101001001001" => q_unbuf <= my_rom(2633);
      when "0101001001010" => q_unbuf <= my_rom(2634);
      when "0101001001011" => q_unbuf <= my_rom(2635);
      when "0101001001100" => q_unbuf <= my_rom(2636);
      when "0101001001101" => q_unbuf <= my_rom(2637);
      when "0101001001110" => q_unbuf <= my_rom(2638);
      when "0101001001111" => q_unbuf <= my_rom(2639);
      when "0101001010000" => q_unbuf <= my_rom(2640);
      when "0101001010001" => q_unbuf <= my_rom(2641);
      when "0101001010010" => q_unbuf <= my_rom(2642);
      when "0101001010011" => q_unbuf <= my_rom(2643);
      when "0101001010100" => q_unbuf <= my_rom(2644);
      when "0101001010101" => q_unbuf <= my_rom(2645);
      when "0101001010110" => q_unbuf <= my_rom(2646);
      when "0101001010111" => q_unbuf <= my_rom(2647);
      when "0101001011000" => q_unbuf <= my_rom(2648);
      when "0101001011001" => q_unbuf <= my_rom(2649);
      when "0101001011010" => q_unbuf <= my_rom(2650);
      when "0101001011011" => q_unbuf <= my_rom(2651);
      when "0101001011100" => q_unbuf <= my_rom(2652);
      when "0101001011101" => q_unbuf <= my_rom(2653);
      when "0101001011110" => q_unbuf <= my_rom(2654);
      when "0101001011111" => q_unbuf <= my_rom(2655);
      when "0101001100000" => q_unbuf <= my_rom(2656);
      when "0101001100001" => q_unbuf <= my_rom(2657);
      when "0101001100010" => q_unbuf <= my_rom(2658);
      when "0101001100011" => q_unbuf <= my_rom(2659);
      when "0101001100100" => q_unbuf <= my_rom(2660);
      when "0101001100101" => q_unbuf <= my_rom(2661);
      when "0101001100110" => q_unbuf <= my_rom(2662);
      when "0101001100111" => q_unbuf <= my_rom(2663);
      when "0101001101000" => q_unbuf <= my_rom(2664);
      when "0101001101001" => q_unbuf <= my_rom(2665);
      when "0101001101010" => q_unbuf <= my_rom(2666);
      when "0101001101011" => q_unbuf <= my_rom(2667);
      when "0101001101100" => q_unbuf <= my_rom(2668);
      when "0101001101101" => q_unbuf <= my_rom(2669);
      when "0101001101110" => q_unbuf <= my_rom(2670);
      when "0101001101111" => q_unbuf <= my_rom(2671);
      when "0101001110000" => q_unbuf <= my_rom(2672);
      when "0101001110001" => q_unbuf <= my_rom(2673);
      when "0101001110010" => q_unbuf <= my_rom(2674);
      when "0101001110011" => q_unbuf <= my_rom(2675);
      when "0101001110100" => q_unbuf <= my_rom(2676);
      when "0101001110101" => q_unbuf <= my_rom(2677);
      when "0101001110110" => q_unbuf <= my_rom(2678);
      when "0101001110111" => q_unbuf <= my_rom(2679);
      when "0101001111000" => q_unbuf <= my_rom(2680);
      when "0101001111001" => q_unbuf <= my_rom(2681);
      when "0101001111010" => q_unbuf <= my_rom(2682);
      when "0101001111011" => q_unbuf <= my_rom(2683);
      when "0101001111100" => q_unbuf <= my_rom(2684);
      when "0101001111101" => q_unbuf <= my_rom(2685);
      when "0101001111110" => q_unbuf <= my_rom(2686);
      when "0101001111111" => q_unbuf <= my_rom(2687);
      when "0101010000000" => q_unbuf <= my_rom(2688);
      when "0101010000001" => q_unbuf <= my_rom(2689);
      when "0101010000010" => q_unbuf <= my_rom(2690);
      when "0101010000011" => q_unbuf <= my_rom(2691);
      when "0101010000100" => q_unbuf <= my_rom(2692);
      when "0101010000101" => q_unbuf <= my_rom(2693);
      when "0101010000110" => q_unbuf <= my_rom(2694);
      when "0101010000111" => q_unbuf <= my_rom(2695);
      when "0101010001000" => q_unbuf <= my_rom(2696);
      when "0101010001001" => q_unbuf <= my_rom(2697);
      when "0101010001010" => q_unbuf <= my_rom(2698);
      when "0101010001011" => q_unbuf <= my_rom(2699);
      when "0101010001100" => q_unbuf <= my_rom(2700);
      when "0101010001101" => q_unbuf <= my_rom(2701);
      when "0101010001110" => q_unbuf <= my_rom(2702);
      when "0101010001111" => q_unbuf <= my_rom(2703);
      when "0101010010000" => q_unbuf <= my_rom(2704);
      when "0101010010001" => q_unbuf <= my_rom(2705);
      when "0101010010010" => q_unbuf <= my_rom(2706);
      when "0101010010011" => q_unbuf <= my_rom(2707);
      when "0101010010100" => q_unbuf <= my_rom(2708);
      when "0101010010101" => q_unbuf <= my_rom(2709);
      when "0101010010110" => q_unbuf <= my_rom(2710);
      when "0101010010111" => q_unbuf <= my_rom(2711);
      when "0101010011000" => q_unbuf <= my_rom(2712);
      when "0101010011001" => q_unbuf <= my_rom(2713);
      when "0101010011010" => q_unbuf <= my_rom(2714);
      when "0101010011011" => q_unbuf <= my_rom(2715);
      when "0101010011100" => q_unbuf <= my_rom(2716);
      when "0101010011101" => q_unbuf <= my_rom(2717);
      when "0101010011110" => q_unbuf <= my_rom(2718);
      when "0101010011111" => q_unbuf <= my_rom(2719);
      when "0101010100000" => q_unbuf <= my_rom(2720);
      when "0101010100001" => q_unbuf <= my_rom(2721);
      when "0101010100010" => q_unbuf <= my_rom(2722);
      when "0101010100011" => q_unbuf <= my_rom(2723);
      when "0101010100100" => q_unbuf <= my_rom(2724);
      when "0101010100101" => q_unbuf <= my_rom(2725);
      when "0101010100110" => q_unbuf <= my_rom(2726);
      when "0101010100111" => q_unbuf <= my_rom(2727);
      when "0101010101000" => q_unbuf <= my_rom(2728);
      when "0101010101001" => q_unbuf <= my_rom(2729);
      when "0101010101010" => q_unbuf <= my_rom(2730);
      when "0101010101011" => q_unbuf <= my_rom(2731);
      when "0101010101100" => q_unbuf <= my_rom(2732);
      when "0101010101101" => q_unbuf <= my_rom(2733);
      when "0101010101110" => q_unbuf <= my_rom(2734);
      when "0101010101111" => q_unbuf <= my_rom(2735);
      when "0101010110000" => q_unbuf <= my_rom(2736);
      when "0101010110001" => q_unbuf <= my_rom(2737);
      when "0101010110010" => q_unbuf <= my_rom(2738);
      when "0101010110011" => q_unbuf <= my_rom(2739);
      when "0101010110100" => q_unbuf <= my_rom(2740);
      when "0101010110101" => q_unbuf <= my_rom(2741);
      when "0101010110110" => q_unbuf <= my_rom(2742);
      when "0101010110111" => q_unbuf <= my_rom(2743);
      when "0101010111000" => q_unbuf <= my_rom(2744);
      when "0101010111001" => q_unbuf <= my_rom(2745);
      when "0101010111010" => q_unbuf <= my_rom(2746);
      when "0101010111011" => q_unbuf <= my_rom(2747);
      when "0101010111100" => q_unbuf <= my_rom(2748);
      when "0101010111101" => q_unbuf <= my_rom(2749);
      when "0101010111110" => q_unbuf <= my_rom(2750);
      when "0101010111111" => q_unbuf <= my_rom(2751);
      when "0101011000000" => q_unbuf <= my_rom(2752);
      when "0101011000001" => q_unbuf <= my_rom(2753);
      when "0101011000010" => q_unbuf <= my_rom(2754);
      when "0101011000011" => q_unbuf <= my_rom(2755);
      when "0101011000100" => q_unbuf <= my_rom(2756);
      when "0101011000101" => q_unbuf <= my_rom(2757);
      when "0101011000110" => q_unbuf <= my_rom(2758);
      when "0101011000111" => q_unbuf <= my_rom(2759);
      when "0101011001000" => q_unbuf <= my_rom(2760);
      when "0101011001001" => q_unbuf <= my_rom(2761);
      when "0101011001010" => q_unbuf <= my_rom(2762);
      when "0101011001011" => q_unbuf <= my_rom(2763);
      when "0101011001100" => q_unbuf <= my_rom(2764);
      when "0101011001101" => q_unbuf <= my_rom(2765);
      when "0101011001110" => q_unbuf <= my_rom(2766);
      when "0101011001111" => q_unbuf <= my_rom(2767);
      when "0101011010000" => q_unbuf <= my_rom(2768);
      when "0101011010001" => q_unbuf <= my_rom(2769);
      when "0101011010010" => q_unbuf <= my_rom(2770);
      when "0101011010011" => q_unbuf <= my_rom(2771);
      when "0101011010100" => q_unbuf <= my_rom(2772);
      when "0101011010101" => q_unbuf <= my_rom(2773);
      when "0101011010110" => q_unbuf <= my_rom(2774);
      when "0101011010111" => q_unbuf <= my_rom(2775);
      when "0101011011000" => q_unbuf <= my_rom(2776);
      when "0101011011001" => q_unbuf <= my_rom(2777);
      when "0101011011010" => q_unbuf <= my_rom(2778);
      when "0101011011011" => q_unbuf <= my_rom(2779);
      when "0101011011100" => q_unbuf <= my_rom(2780);
      when "0101011011101" => q_unbuf <= my_rom(2781);
      when "0101011011110" => q_unbuf <= my_rom(2782);
      when "0101011011111" => q_unbuf <= my_rom(2783);
      when "0101011100000" => q_unbuf <= my_rom(2784);
      when "0101011100001" => q_unbuf <= my_rom(2785);
      when "0101011100010" => q_unbuf <= my_rom(2786);
      when "0101011100011" => q_unbuf <= my_rom(2787);
      when "0101011100100" => q_unbuf <= my_rom(2788);
      when "0101011100101" => q_unbuf <= my_rom(2789);
      when "0101011100110" => q_unbuf <= my_rom(2790);
      when "0101011100111" => q_unbuf <= my_rom(2791);
      when "0101011101000" => q_unbuf <= my_rom(2792);
      when "0101011101001" => q_unbuf <= my_rom(2793);
      when "0101011101010" => q_unbuf <= my_rom(2794);
      when "0101011101011" => q_unbuf <= my_rom(2795);
      when "0101011101100" => q_unbuf <= my_rom(2796);
      when "0101011101101" => q_unbuf <= my_rom(2797);
      when "0101011101110" => q_unbuf <= my_rom(2798);
      when "0101011101111" => q_unbuf <= my_rom(2799);
      when "0101011110000" => q_unbuf <= my_rom(2800);
      when "0101011110001" => q_unbuf <= my_rom(2801);
      when "0101011110010" => q_unbuf <= my_rom(2802);
      when "0101011110011" => q_unbuf <= my_rom(2803);
      when "0101011110100" => q_unbuf <= my_rom(2804);
      when "0101011110101" => q_unbuf <= my_rom(2805);
      when "0101011110110" => q_unbuf <= my_rom(2806);
      when "0101011110111" => q_unbuf <= my_rom(2807);
      when "0101011111000" => q_unbuf <= my_rom(2808);
      when "0101011111001" => q_unbuf <= my_rom(2809);
      when "0101011111010" => q_unbuf <= my_rom(2810);
      when "0101011111011" => q_unbuf <= my_rom(2811);
      when "0101011111100" => q_unbuf <= my_rom(2812);
      when "0101011111101" => q_unbuf <= my_rom(2813);
      when "0101011111110" => q_unbuf <= my_rom(2814);
      when "0101011111111" => q_unbuf <= my_rom(2815);
      when "0101100000000" => q_unbuf <= my_rom(2816);
      when "0101100000001" => q_unbuf <= my_rom(2817);
      when "0101100000010" => q_unbuf <= my_rom(2818);
      when "0101100000011" => q_unbuf <= my_rom(2819);
      when "0101100000100" => q_unbuf <= my_rom(2820);
      when "0101100000101" => q_unbuf <= my_rom(2821);
      when "0101100000110" => q_unbuf <= my_rom(2822);
      when "0101100000111" => q_unbuf <= my_rom(2823);
      when "0101100001000" => q_unbuf <= my_rom(2824);
      when "0101100001001" => q_unbuf <= my_rom(2825);
      when "0101100001010" => q_unbuf <= my_rom(2826);
      when "0101100001011" => q_unbuf <= my_rom(2827);
      when "0101100001100" => q_unbuf <= my_rom(2828);
      when "0101100001101" => q_unbuf <= my_rom(2829);
      when "0101100001110" => q_unbuf <= my_rom(2830);
      when "0101100001111" => q_unbuf <= my_rom(2831);
      when "0101100010000" => q_unbuf <= my_rom(2832);
      when "0101100010001" => q_unbuf <= my_rom(2833);
      when "0101100010010" => q_unbuf <= my_rom(2834);
      when "0101100010011" => q_unbuf <= my_rom(2835);
      when "0101100010100" => q_unbuf <= my_rom(2836);
      when "0101100010101" => q_unbuf <= my_rom(2837);
      when "0101100010110" => q_unbuf <= my_rom(2838);
      when "0101100010111" => q_unbuf <= my_rom(2839);
      when "0101100011000" => q_unbuf <= my_rom(2840);
      when "0101100011001" => q_unbuf <= my_rom(2841);
      when "0101100011010" => q_unbuf <= my_rom(2842);
      when "0101100011011" => q_unbuf <= my_rom(2843);
      when "0101100011100" => q_unbuf <= my_rom(2844);
      when "0101100011101" => q_unbuf <= my_rom(2845);
      when "0101100011110" => q_unbuf <= my_rom(2846);
      when "0101100011111" => q_unbuf <= my_rom(2847);
      when "0101100100000" => q_unbuf <= my_rom(2848);
      when "0101100100001" => q_unbuf <= my_rom(2849);
      when "0101100100010" => q_unbuf <= my_rom(2850);
      when "0101100100011" => q_unbuf <= my_rom(2851);
      when "0101100100100" => q_unbuf <= my_rom(2852);
      when "0101100100101" => q_unbuf <= my_rom(2853);
      when "0101100100110" => q_unbuf <= my_rom(2854);
      when "0101100100111" => q_unbuf <= my_rom(2855);
      when "0101100101000" => q_unbuf <= my_rom(2856);
      when "0101100101001" => q_unbuf <= my_rom(2857);
      when "0101100101010" => q_unbuf <= my_rom(2858);
      when "0101100101011" => q_unbuf <= my_rom(2859);
      when "0101100101100" => q_unbuf <= my_rom(2860);
      when "0101100101101" => q_unbuf <= my_rom(2861);
      when "0101100101110" => q_unbuf <= my_rom(2862);
      when "0101100101111" => q_unbuf <= my_rom(2863);
      when "0101100110000" => q_unbuf <= my_rom(2864);
      when "0101100110001" => q_unbuf <= my_rom(2865);
      when "0101100110010" => q_unbuf <= my_rom(2866);
      when "0101100110011" => q_unbuf <= my_rom(2867);
      when "0101100110100" => q_unbuf <= my_rom(2868);
      when "0101100110101" => q_unbuf <= my_rom(2869);
      when "0101100110110" => q_unbuf <= my_rom(2870);
      when "0101100110111" => q_unbuf <= my_rom(2871);
      when "0101100111000" => q_unbuf <= my_rom(2872);
      when "0101100111001" => q_unbuf <= my_rom(2873);
      when "0101100111010" => q_unbuf <= my_rom(2874);
      when "0101100111011" => q_unbuf <= my_rom(2875);
      when "0101100111100" => q_unbuf <= my_rom(2876);
      when "0101100111101" => q_unbuf <= my_rom(2877);
      when "0101100111110" => q_unbuf <= my_rom(2878);
      when "0101100111111" => q_unbuf <= my_rom(2879);
      when "0101101000000" => q_unbuf <= my_rom(2880);
      when "0101101000001" => q_unbuf <= my_rom(2881);
      when "0101101000010" => q_unbuf <= my_rom(2882);
      when "0101101000011" => q_unbuf <= my_rom(2883);
      when "0101101000100" => q_unbuf <= my_rom(2884);
      when "0101101000101" => q_unbuf <= my_rom(2885);
      when "0101101000110" => q_unbuf <= my_rom(2886);
      when "0101101000111" => q_unbuf <= my_rom(2887);
      when "0101101001000" => q_unbuf <= my_rom(2888);
      when "0101101001001" => q_unbuf <= my_rom(2889);
      when "0101101001010" => q_unbuf <= my_rom(2890);
      when "0101101001011" => q_unbuf <= my_rom(2891);
      when "0101101001100" => q_unbuf <= my_rom(2892);
      when "0101101001101" => q_unbuf <= my_rom(2893);
      when "0101101001110" => q_unbuf <= my_rom(2894);
      when "0101101001111" => q_unbuf <= my_rom(2895);
      when "0101101010000" => q_unbuf <= my_rom(2896);
      when "0101101010001" => q_unbuf <= my_rom(2897);
      when "0101101010010" => q_unbuf <= my_rom(2898);
      when "0101101010011" => q_unbuf <= my_rom(2899);
      when "0101101010100" => q_unbuf <= my_rom(2900);
      when "0101101010101" => q_unbuf <= my_rom(2901);
      when "0101101010110" => q_unbuf <= my_rom(2902);
      when "0101101010111" => q_unbuf <= my_rom(2903);
      when "0101101011000" => q_unbuf <= my_rom(2904);
      when "0101101011001" => q_unbuf <= my_rom(2905);
      when "0101101011010" => q_unbuf <= my_rom(2906);
      when "0101101011011" => q_unbuf <= my_rom(2907);
      when "0101101011100" => q_unbuf <= my_rom(2908);
      when "0101101011101" => q_unbuf <= my_rom(2909);
      when "0101101011110" => q_unbuf <= my_rom(2910);
      when "0101101011111" => q_unbuf <= my_rom(2911);
      when "0101101100000" => q_unbuf <= my_rom(2912);
      when "0101101100001" => q_unbuf <= my_rom(2913);
      when "0101101100010" => q_unbuf <= my_rom(2914);
      when "0101101100011" => q_unbuf <= my_rom(2915);
      when "0101101100100" => q_unbuf <= my_rom(2916);
      when "0101101100101" => q_unbuf <= my_rom(2917);
      when "0101101100110" => q_unbuf <= my_rom(2918);
      when "0101101100111" => q_unbuf <= my_rom(2919);
      when "0101101101000" => q_unbuf <= my_rom(2920);
      when "0101101101001" => q_unbuf <= my_rom(2921);
      when "0101101101010" => q_unbuf <= my_rom(2922);
      when "0101101101011" => q_unbuf <= my_rom(2923);
      when "0101101101100" => q_unbuf <= my_rom(2924);
      when "0101101101101" => q_unbuf <= my_rom(2925);
      when "0101101101110" => q_unbuf <= my_rom(2926);
      when "0101101101111" => q_unbuf <= my_rom(2927);
      when "0101101110000" => q_unbuf <= my_rom(2928);
      when "0101101110001" => q_unbuf <= my_rom(2929);
      when "0101101110010" => q_unbuf <= my_rom(2930);
      when "0101101110011" => q_unbuf <= my_rom(2931);
      when "0101101110100" => q_unbuf <= my_rom(2932);
      when "0101101110101" => q_unbuf <= my_rom(2933);
      when "0101101110110" => q_unbuf <= my_rom(2934);
      when "0101101110111" => q_unbuf <= my_rom(2935);
      when "0101101111000" => q_unbuf <= my_rom(2936);
      when "0101101111001" => q_unbuf <= my_rom(2937);
      when "0101101111010" => q_unbuf <= my_rom(2938);
      when "0101101111011" => q_unbuf <= my_rom(2939);
      when "0101101111100" => q_unbuf <= my_rom(2940);
      when "0101101111101" => q_unbuf <= my_rom(2941);
      when "0101101111110" => q_unbuf <= my_rom(2942);
      when "0101101111111" => q_unbuf <= my_rom(2943);
      when "0101110000000" => q_unbuf <= my_rom(2944);
      when "0101110000001" => q_unbuf <= my_rom(2945);
      when "0101110000010" => q_unbuf <= my_rom(2946);
      when "0101110000011" => q_unbuf <= my_rom(2947);
      when "0101110000100" => q_unbuf <= my_rom(2948);
      when "0101110000101" => q_unbuf <= my_rom(2949);
      when "0101110000110" => q_unbuf <= my_rom(2950);
      when "0101110000111" => q_unbuf <= my_rom(2951);
      when "0101110001000" => q_unbuf <= my_rom(2952);
      when "0101110001001" => q_unbuf <= my_rom(2953);
      when "0101110001010" => q_unbuf <= my_rom(2954);
      when "0101110001011" => q_unbuf <= my_rom(2955);
      when "0101110001100" => q_unbuf <= my_rom(2956);
      when "0101110001101" => q_unbuf <= my_rom(2957);
      when "0101110001110" => q_unbuf <= my_rom(2958);
      when "0101110001111" => q_unbuf <= my_rom(2959);
      when "0101110010000" => q_unbuf <= my_rom(2960);
      when "0101110010001" => q_unbuf <= my_rom(2961);
      when "0101110010010" => q_unbuf <= my_rom(2962);
      when "0101110010011" => q_unbuf <= my_rom(2963);
      when "0101110010100" => q_unbuf <= my_rom(2964);
      when "0101110010101" => q_unbuf <= my_rom(2965);
      when "0101110010110" => q_unbuf <= my_rom(2966);
      when "0101110010111" => q_unbuf <= my_rom(2967);
      when "0101110011000" => q_unbuf <= my_rom(2968);
      when "0101110011001" => q_unbuf <= my_rom(2969);
      when "0101110011010" => q_unbuf <= my_rom(2970);
      when "0101110011011" => q_unbuf <= my_rom(2971);
      when "0101110011100" => q_unbuf <= my_rom(2972);
      when "0101110011101" => q_unbuf <= my_rom(2973);
      when "0101110011110" => q_unbuf <= my_rom(2974);
      when "0101110011111" => q_unbuf <= my_rom(2975);
      when "0101110100000" => q_unbuf <= my_rom(2976);
      when "0101110100001" => q_unbuf <= my_rom(2977);
      when "0101110100010" => q_unbuf <= my_rom(2978);
      when "0101110100011" => q_unbuf <= my_rom(2979);
      when "0101110100100" => q_unbuf <= my_rom(2980);
      when "0101110100101" => q_unbuf <= my_rom(2981);
      when "0101110100110" => q_unbuf <= my_rom(2982);
      when "0101110100111" => q_unbuf <= my_rom(2983);
      when "0101110101000" => q_unbuf <= my_rom(2984);
      when "0101110101001" => q_unbuf <= my_rom(2985);
      when "0101110101010" => q_unbuf <= my_rom(2986);
      when "0101110101011" => q_unbuf <= my_rom(2987);
      when "0101110101100" => q_unbuf <= my_rom(2988);
      when "0101110101101" => q_unbuf <= my_rom(2989);
      when "0101110101110" => q_unbuf <= my_rom(2990);
      when "0101110101111" => q_unbuf <= my_rom(2991);
      when "0101110110000" => q_unbuf <= my_rom(2992);
      when "0101110110001" => q_unbuf <= my_rom(2993);
      when "0101110110010" => q_unbuf <= my_rom(2994);
      when "0101110110011" => q_unbuf <= my_rom(2995);
      when "0101110110100" => q_unbuf <= my_rom(2996);
      when "0101110110101" => q_unbuf <= my_rom(2997);
      when "0101110110110" => q_unbuf <= my_rom(2998);
      when "0101110110111" => q_unbuf <= my_rom(2999);
      when "0101110111000" => q_unbuf <= my_rom(3000);
      when "0101110111001" => q_unbuf <= my_rom(3001);
      when "0101110111010" => q_unbuf <= my_rom(3002);
      when "0101110111011" => q_unbuf <= my_rom(3003);
      when "0101110111100" => q_unbuf <= my_rom(3004);
      when "0101110111101" => q_unbuf <= my_rom(3005);
      when "0101110111110" => q_unbuf <= my_rom(3006);
      when "0101110111111" => q_unbuf <= my_rom(3007);
      when "0101111000000" => q_unbuf <= my_rom(3008);
      when "0101111000001" => q_unbuf <= my_rom(3009);
      when "0101111000010" => q_unbuf <= my_rom(3010);
      when "0101111000011" => q_unbuf <= my_rom(3011);
      when "0101111000100" => q_unbuf <= my_rom(3012);
      when "0101111000101" => q_unbuf <= my_rom(3013);
      when "0101111000110" => q_unbuf <= my_rom(3014);
      when "0101111000111" => q_unbuf <= my_rom(3015);
      when "0101111001000" => q_unbuf <= my_rom(3016);
      when "0101111001001" => q_unbuf <= my_rom(3017);
      when "0101111001010" => q_unbuf <= my_rom(3018);
      when "0101111001011" => q_unbuf <= my_rom(3019);
      when "0101111001100" => q_unbuf <= my_rom(3020);
      when "0101111001101" => q_unbuf <= my_rom(3021);
      when "0101111001110" => q_unbuf <= my_rom(3022);
      when "0101111001111" => q_unbuf <= my_rom(3023);
      when "0101111010000" => q_unbuf <= my_rom(3024);
      when "0101111010001" => q_unbuf <= my_rom(3025);
      when "0101111010010" => q_unbuf <= my_rom(3026);
      when "0101111010011" => q_unbuf <= my_rom(3027);
      when "0101111010100" => q_unbuf <= my_rom(3028);
      when "0101111010101" => q_unbuf <= my_rom(3029);
      when "0101111010110" => q_unbuf <= my_rom(3030);
      when "0101111010111" => q_unbuf <= my_rom(3031);
      when "0101111011000" => q_unbuf <= my_rom(3032);
      when "0101111011001" => q_unbuf <= my_rom(3033);
      when "0101111011010" => q_unbuf <= my_rom(3034);
      when "0101111011011" => q_unbuf <= my_rom(3035);
      when "0101111011100" => q_unbuf <= my_rom(3036);
      when "0101111011101" => q_unbuf <= my_rom(3037);
      when "0101111011110" => q_unbuf <= my_rom(3038);
      when "0101111011111" => q_unbuf <= my_rom(3039);
      when "0101111100000" => q_unbuf <= my_rom(3040);
      when "0101111100001" => q_unbuf <= my_rom(3041);
      when "0101111100010" => q_unbuf <= my_rom(3042);
      when "0101111100011" => q_unbuf <= my_rom(3043);
      when "0101111100100" => q_unbuf <= my_rom(3044);
      when "0101111100101" => q_unbuf <= my_rom(3045);
      when "0101111100110" => q_unbuf <= my_rom(3046);
      when "0101111100111" => q_unbuf <= my_rom(3047);
      when "0101111101000" => q_unbuf <= my_rom(3048);
      when "0101111101001" => q_unbuf <= my_rom(3049);
      when "0101111101010" => q_unbuf <= my_rom(3050);
      when "0101111101011" => q_unbuf <= my_rom(3051);
      when "0101111101100" => q_unbuf <= my_rom(3052);
      when "0101111101101" => q_unbuf <= my_rom(3053);
      when "0101111101110" => q_unbuf <= my_rom(3054);
      when "0101111101111" => q_unbuf <= my_rom(3055);
      when "0101111110000" => q_unbuf <= my_rom(3056);
      when "0101111110001" => q_unbuf <= my_rom(3057);
      when "0101111110010" => q_unbuf <= my_rom(3058);
      when "0101111110011" => q_unbuf <= my_rom(3059);
      when "0101111110100" => q_unbuf <= my_rom(3060);
      when "0101111110101" => q_unbuf <= my_rom(3061);
      when "0101111110110" => q_unbuf <= my_rom(3062);
      when "0101111110111" => q_unbuf <= my_rom(3063);
      when "0101111111000" => q_unbuf <= my_rom(3064);
      when "0101111111001" => q_unbuf <= my_rom(3065);
      when "0101111111010" => q_unbuf <= my_rom(3066);
      when "0101111111011" => q_unbuf <= my_rom(3067);
      when "0101111111100" => q_unbuf <= my_rom(3068);
      when "0101111111101" => q_unbuf <= my_rom(3069);
      when "0101111111110" => q_unbuf <= my_rom(3070);
      when "0101111111111" => q_unbuf <= my_rom(3071);
      when "0110000000000" => q_unbuf <= my_rom(3072);
      when "0110000000001" => q_unbuf <= my_rom(3073);
      when "0110000000010" => q_unbuf <= my_rom(3074);
      when "0110000000011" => q_unbuf <= my_rom(3075);
      when "0110000000100" => q_unbuf <= my_rom(3076);
      when "0110000000101" => q_unbuf <= my_rom(3077);
      when "0110000000110" => q_unbuf <= my_rom(3078);
      when "0110000000111" => q_unbuf <= my_rom(3079);
      when "0110000001000" => q_unbuf <= my_rom(3080);
      when "0110000001001" => q_unbuf <= my_rom(3081);
      when "0110000001010" => q_unbuf <= my_rom(3082);
      when "0110000001011" => q_unbuf <= my_rom(3083);
      when "0110000001100" => q_unbuf <= my_rom(3084);
      when "0110000001101" => q_unbuf <= my_rom(3085);
      when "0110000001110" => q_unbuf <= my_rom(3086);
      when "0110000001111" => q_unbuf <= my_rom(3087);
      when "0110000010000" => q_unbuf <= my_rom(3088);
      when "0110000010001" => q_unbuf <= my_rom(3089);
      when "0110000010010" => q_unbuf <= my_rom(3090);
      when "0110000010011" => q_unbuf <= my_rom(3091);
      when "0110000010100" => q_unbuf <= my_rom(3092);
      when "0110000010101" => q_unbuf <= my_rom(3093);
      when "0110000010110" => q_unbuf <= my_rom(3094);
      when "0110000010111" => q_unbuf <= my_rom(3095);
      when "0110000011000" => q_unbuf <= my_rom(3096);
      when "0110000011001" => q_unbuf <= my_rom(3097);
      when "0110000011010" => q_unbuf <= my_rom(3098);
      when "0110000011011" => q_unbuf <= my_rom(3099);
      when "0110000011100" => q_unbuf <= my_rom(3100);
      when "0110000011101" => q_unbuf <= my_rom(3101);
      when "0110000011110" => q_unbuf <= my_rom(3102);
      when "0110000011111" => q_unbuf <= my_rom(3103);
      when "0110000100000" => q_unbuf <= my_rom(3104);
      when "0110000100001" => q_unbuf <= my_rom(3105);
      when "0110000100010" => q_unbuf <= my_rom(3106);
      when "0110000100011" => q_unbuf <= my_rom(3107);
      when "0110000100100" => q_unbuf <= my_rom(3108);
      when "0110000100101" => q_unbuf <= my_rom(3109);
      when "0110000100110" => q_unbuf <= my_rom(3110);
      when "0110000100111" => q_unbuf <= my_rom(3111);
      when "0110000101000" => q_unbuf <= my_rom(3112);
      when "0110000101001" => q_unbuf <= my_rom(3113);
      when "0110000101010" => q_unbuf <= my_rom(3114);
      when "0110000101011" => q_unbuf <= my_rom(3115);
      when "0110000101100" => q_unbuf <= my_rom(3116);
      when "0110000101101" => q_unbuf <= my_rom(3117);
      when "0110000101110" => q_unbuf <= my_rom(3118);
      when "0110000101111" => q_unbuf <= my_rom(3119);
      when "0110000110000" => q_unbuf <= my_rom(3120);
      when "0110000110001" => q_unbuf <= my_rom(3121);
      when "0110000110010" => q_unbuf <= my_rom(3122);
      when "0110000110011" => q_unbuf <= my_rom(3123);
      when "0110000110100" => q_unbuf <= my_rom(3124);
      when "0110000110101" => q_unbuf <= my_rom(3125);
      when "0110000110110" => q_unbuf <= my_rom(3126);
      when "0110000110111" => q_unbuf <= my_rom(3127);
      when "0110000111000" => q_unbuf <= my_rom(3128);
      when "0110000111001" => q_unbuf <= my_rom(3129);
      when "0110000111010" => q_unbuf <= my_rom(3130);
      when "0110000111011" => q_unbuf <= my_rom(3131);
      when "0110000111100" => q_unbuf <= my_rom(3132);
      when "0110000111101" => q_unbuf <= my_rom(3133);
      when "0110000111110" => q_unbuf <= my_rom(3134);
      when "0110000111111" => q_unbuf <= my_rom(3135);
      when "0110001000000" => q_unbuf <= my_rom(3136);
      when "0110001000001" => q_unbuf <= my_rom(3137);
      when "0110001000010" => q_unbuf <= my_rom(3138);
      when "0110001000011" => q_unbuf <= my_rom(3139);
      when "0110001000100" => q_unbuf <= my_rom(3140);
      when "0110001000101" => q_unbuf <= my_rom(3141);
      when "0110001000110" => q_unbuf <= my_rom(3142);
      when "0110001000111" => q_unbuf <= my_rom(3143);
      when "0110001001000" => q_unbuf <= my_rom(3144);
      when "0110001001001" => q_unbuf <= my_rom(3145);
      when "0110001001010" => q_unbuf <= my_rom(3146);
      when "0110001001011" => q_unbuf <= my_rom(3147);
      when "0110001001100" => q_unbuf <= my_rom(3148);
      when "0110001001101" => q_unbuf <= my_rom(3149);
      when "0110001001110" => q_unbuf <= my_rom(3150);
      when "0110001001111" => q_unbuf <= my_rom(3151);
      when "0110001010000" => q_unbuf <= my_rom(3152);
      when "0110001010001" => q_unbuf <= my_rom(3153);
      when "0110001010010" => q_unbuf <= my_rom(3154);
      when "0110001010011" => q_unbuf <= my_rom(3155);
      when "0110001010100" => q_unbuf <= my_rom(3156);
      when "0110001010101" => q_unbuf <= my_rom(3157);
      when "0110001010110" => q_unbuf <= my_rom(3158);
      when "0110001010111" => q_unbuf <= my_rom(3159);
      when "0110001011000" => q_unbuf <= my_rom(3160);
      when "0110001011001" => q_unbuf <= my_rom(3161);
      when "0110001011010" => q_unbuf <= my_rom(3162);
      when "0110001011011" => q_unbuf <= my_rom(3163);
      when "0110001011100" => q_unbuf <= my_rom(3164);
      when "0110001011101" => q_unbuf <= my_rom(3165);
      when "0110001011110" => q_unbuf <= my_rom(3166);
      when "0110001011111" => q_unbuf <= my_rom(3167);
      when "0110001100000" => q_unbuf <= my_rom(3168);
      when "0110001100001" => q_unbuf <= my_rom(3169);
      when "0110001100010" => q_unbuf <= my_rom(3170);
      when "0110001100011" => q_unbuf <= my_rom(3171);
      when "0110001100100" => q_unbuf <= my_rom(3172);
      when "0110001100101" => q_unbuf <= my_rom(3173);
      when "0110001100110" => q_unbuf <= my_rom(3174);
      when "0110001100111" => q_unbuf <= my_rom(3175);
      when "0110001101000" => q_unbuf <= my_rom(3176);
      when "0110001101001" => q_unbuf <= my_rom(3177);
      when "0110001101010" => q_unbuf <= my_rom(3178);
      when "0110001101011" => q_unbuf <= my_rom(3179);
      when "0110001101100" => q_unbuf <= my_rom(3180);
      when "0110001101101" => q_unbuf <= my_rom(3181);
      when "0110001101110" => q_unbuf <= my_rom(3182);
      when "0110001101111" => q_unbuf <= my_rom(3183);
      when "0110001110000" => q_unbuf <= my_rom(3184);
      when "0110001110001" => q_unbuf <= my_rom(3185);
      when "0110001110010" => q_unbuf <= my_rom(3186);
      when "0110001110011" => q_unbuf <= my_rom(3187);
      when "0110001110100" => q_unbuf <= my_rom(3188);
      when "0110001110101" => q_unbuf <= my_rom(3189);
      when "0110001110110" => q_unbuf <= my_rom(3190);
      when "0110001110111" => q_unbuf <= my_rom(3191);
      when "0110001111000" => q_unbuf <= my_rom(3192);
      when "0110001111001" => q_unbuf <= my_rom(3193);
      when "0110001111010" => q_unbuf <= my_rom(3194);
      when "0110001111011" => q_unbuf <= my_rom(3195);
      when "0110001111100" => q_unbuf <= my_rom(3196);
      when "0110001111101" => q_unbuf <= my_rom(3197);
      when "0110001111110" => q_unbuf <= my_rom(3198);
      when "0110001111111" => q_unbuf <= my_rom(3199);
      when "0110010000000" => q_unbuf <= my_rom(3200);
      when "0110010000001" => q_unbuf <= my_rom(3201);
      when "0110010000010" => q_unbuf <= my_rom(3202);
      when "0110010000011" => q_unbuf <= my_rom(3203);
      when "0110010000100" => q_unbuf <= my_rom(3204);
      when "0110010000101" => q_unbuf <= my_rom(3205);
      when "0110010000110" => q_unbuf <= my_rom(3206);
      when "0110010000111" => q_unbuf <= my_rom(3207);
      when "0110010001000" => q_unbuf <= my_rom(3208);
      when "0110010001001" => q_unbuf <= my_rom(3209);
      when "0110010001010" => q_unbuf <= my_rom(3210);
      when "0110010001011" => q_unbuf <= my_rom(3211);
      when "0110010001100" => q_unbuf <= my_rom(3212);
      when "0110010001101" => q_unbuf <= my_rom(3213);
      when "0110010001110" => q_unbuf <= my_rom(3214);
      when "0110010001111" => q_unbuf <= my_rom(3215);
      when "0110010010000" => q_unbuf <= my_rom(3216);
      when "0110010010001" => q_unbuf <= my_rom(3217);
      when "0110010010010" => q_unbuf <= my_rom(3218);
      when "0110010010011" => q_unbuf <= my_rom(3219);
      when "0110010010100" => q_unbuf <= my_rom(3220);
      when "0110010010101" => q_unbuf <= my_rom(3221);
      when "0110010010110" => q_unbuf <= my_rom(3222);
      when "0110010010111" => q_unbuf <= my_rom(3223);
      when "0110010011000" => q_unbuf <= my_rom(3224);
      when "0110010011001" => q_unbuf <= my_rom(3225);
      when "0110010011010" => q_unbuf <= my_rom(3226);
      when "0110010011011" => q_unbuf <= my_rom(3227);
      when "0110010011100" => q_unbuf <= my_rom(3228);
      when "0110010011101" => q_unbuf <= my_rom(3229);
      when "0110010011110" => q_unbuf <= my_rom(3230);
      when "0110010011111" => q_unbuf <= my_rom(3231);
      when "0110010100000" => q_unbuf <= my_rom(3232);
      when "0110010100001" => q_unbuf <= my_rom(3233);
      when "0110010100010" => q_unbuf <= my_rom(3234);
      when "0110010100011" => q_unbuf <= my_rom(3235);
      when "0110010100100" => q_unbuf <= my_rom(3236);
      when "0110010100101" => q_unbuf <= my_rom(3237);
      when "0110010100110" => q_unbuf <= my_rom(3238);
      when "0110010100111" => q_unbuf <= my_rom(3239);
      when "0110010101000" => q_unbuf <= my_rom(3240);
      when "0110010101001" => q_unbuf <= my_rom(3241);
      when "0110010101010" => q_unbuf <= my_rom(3242);
      when "0110010101011" => q_unbuf <= my_rom(3243);
      when "0110010101100" => q_unbuf <= my_rom(3244);
      when "0110010101101" => q_unbuf <= my_rom(3245);
      when "0110010101110" => q_unbuf <= my_rom(3246);
      when "0110010101111" => q_unbuf <= my_rom(3247);
      when "0110010110000" => q_unbuf <= my_rom(3248);
      when "0110010110001" => q_unbuf <= my_rom(3249);
      when "0110010110010" => q_unbuf <= my_rom(3250);
      when "0110010110011" => q_unbuf <= my_rom(3251);
      when "0110010110100" => q_unbuf <= my_rom(3252);
      when "0110010110101" => q_unbuf <= my_rom(3253);
      when "0110010110110" => q_unbuf <= my_rom(3254);
      when "0110010110111" => q_unbuf <= my_rom(3255);
      when "0110010111000" => q_unbuf <= my_rom(3256);
      when "0110010111001" => q_unbuf <= my_rom(3257);
      when "0110010111010" => q_unbuf <= my_rom(3258);
      when "0110010111011" => q_unbuf <= my_rom(3259);
      when "0110010111100" => q_unbuf <= my_rom(3260);
      when "0110010111101" => q_unbuf <= my_rom(3261);
      when "0110010111110" => q_unbuf <= my_rom(3262);
      when "0110010111111" => q_unbuf <= my_rom(3263);
      when "0110011000000" => q_unbuf <= my_rom(3264);
      when "0110011000001" => q_unbuf <= my_rom(3265);
      when "0110011000010" => q_unbuf <= my_rom(3266);
      when "0110011000011" => q_unbuf <= my_rom(3267);
      when "0110011000100" => q_unbuf <= my_rom(3268);
      when "0110011000101" => q_unbuf <= my_rom(3269);
      when "0110011000110" => q_unbuf <= my_rom(3270);
      when "0110011000111" => q_unbuf <= my_rom(3271);
      when "0110011001000" => q_unbuf <= my_rom(3272);
      when "0110011001001" => q_unbuf <= my_rom(3273);
      when "0110011001010" => q_unbuf <= my_rom(3274);
      when "0110011001011" => q_unbuf <= my_rom(3275);
      when "0110011001100" => q_unbuf <= my_rom(3276);
      when "0110011001101" => q_unbuf <= my_rom(3277);
      when "0110011001110" => q_unbuf <= my_rom(3278);
      when "0110011001111" => q_unbuf <= my_rom(3279);
      when "0110011010000" => q_unbuf <= my_rom(3280);
      when "0110011010001" => q_unbuf <= my_rom(3281);
      when "0110011010010" => q_unbuf <= my_rom(3282);
      when "0110011010011" => q_unbuf <= my_rom(3283);
      when "0110011010100" => q_unbuf <= my_rom(3284);
      when "0110011010101" => q_unbuf <= my_rom(3285);
      when "0110011010110" => q_unbuf <= my_rom(3286);
      when "0110011010111" => q_unbuf <= my_rom(3287);
      when "0110011011000" => q_unbuf <= my_rom(3288);
      when "0110011011001" => q_unbuf <= my_rom(3289);
      when "0110011011010" => q_unbuf <= my_rom(3290);
      when "0110011011011" => q_unbuf <= my_rom(3291);
      when "0110011011100" => q_unbuf <= my_rom(3292);
      when "0110011011101" => q_unbuf <= my_rom(3293);
      when "0110011011110" => q_unbuf <= my_rom(3294);
      when "0110011011111" => q_unbuf <= my_rom(3295);
      when "0110011100000" => q_unbuf <= my_rom(3296);
      when "0110011100001" => q_unbuf <= my_rom(3297);
      when "0110011100010" => q_unbuf <= my_rom(3298);
      when "0110011100011" => q_unbuf <= my_rom(3299);
      when "0110011100100" => q_unbuf <= my_rom(3300);
      when "0110011100101" => q_unbuf <= my_rom(3301);
      when "0110011100110" => q_unbuf <= my_rom(3302);
      when "0110011100111" => q_unbuf <= my_rom(3303);
      when "0110011101000" => q_unbuf <= my_rom(3304);
      when "0110011101001" => q_unbuf <= my_rom(3305);
      when "0110011101010" => q_unbuf <= my_rom(3306);
      when "0110011101011" => q_unbuf <= my_rom(3307);
      when "0110011101100" => q_unbuf <= my_rom(3308);
      when "0110011101101" => q_unbuf <= my_rom(3309);
      when "0110011101110" => q_unbuf <= my_rom(3310);
      when "0110011101111" => q_unbuf <= my_rom(3311);
      when "0110011110000" => q_unbuf <= my_rom(3312);
      when "0110011110001" => q_unbuf <= my_rom(3313);
      when "0110011110010" => q_unbuf <= my_rom(3314);
      when "0110011110011" => q_unbuf <= my_rom(3315);
      when "0110011110100" => q_unbuf <= my_rom(3316);
      when "0110011110101" => q_unbuf <= my_rom(3317);
      when "0110011110110" => q_unbuf <= my_rom(3318);
      when "0110011110111" => q_unbuf <= my_rom(3319);
      when "0110011111000" => q_unbuf <= my_rom(3320);
      when "0110011111001" => q_unbuf <= my_rom(3321);
      when "0110011111010" => q_unbuf <= my_rom(3322);
      when "0110011111011" => q_unbuf <= my_rom(3323);
      when "0110011111100" => q_unbuf <= my_rom(3324);
      when "0110011111101" => q_unbuf <= my_rom(3325);
      when "0110011111110" => q_unbuf <= my_rom(3326);
      when "0110011111111" => q_unbuf <= my_rom(3327);
      when "0110100000000" => q_unbuf <= my_rom(3328);
      when "0110100000001" => q_unbuf <= my_rom(3329);
      when "0110100000010" => q_unbuf <= my_rom(3330);
      when "0110100000011" => q_unbuf <= my_rom(3331);
      when "0110100000100" => q_unbuf <= my_rom(3332);
      when "0110100000101" => q_unbuf <= my_rom(3333);
      when "0110100000110" => q_unbuf <= my_rom(3334);
      when "0110100000111" => q_unbuf <= my_rom(3335);
      when "0110100001000" => q_unbuf <= my_rom(3336);
      when "0110100001001" => q_unbuf <= my_rom(3337);
      when "0110100001010" => q_unbuf <= my_rom(3338);
      when "0110100001011" => q_unbuf <= my_rom(3339);
      when "0110100001100" => q_unbuf <= my_rom(3340);
      when "0110100001101" => q_unbuf <= my_rom(3341);
      when "0110100001110" => q_unbuf <= my_rom(3342);
      when "0110100001111" => q_unbuf <= my_rom(3343);
      when "0110100010000" => q_unbuf <= my_rom(3344);
      when "0110100010001" => q_unbuf <= my_rom(3345);
      when "0110100010010" => q_unbuf <= my_rom(3346);
      when "0110100010011" => q_unbuf <= my_rom(3347);
      when "0110100010100" => q_unbuf <= my_rom(3348);
      when "0110100010101" => q_unbuf <= my_rom(3349);
      when "0110100010110" => q_unbuf <= my_rom(3350);
      when "0110100010111" => q_unbuf <= my_rom(3351);
      when "0110100011000" => q_unbuf <= my_rom(3352);
      when "0110100011001" => q_unbuf <= my_rom(3353);
      when "0110100011010" => q_unbuf <= my_rom(3354);
      when "0110100011011" => q_unbuf <= my_rom(3355);
      when "0110100011100" => q_unbuf <= my_rom(3356);
      when "0110100011101" => q_unbuf <= my_rom(3357);
      when "0110100011110" => q_unbuf <= my_rom(3358);
      when "0110100011111" => q_unbuf <= my_rom(3359);
      when "0110100100000" => q_unbuf <= my_rom(3360);
      when "0110100100001" => q_unbuf <= my_rom(3361);
      when "0110100100010" => q_unbuf <= my_rom(3362);
      when "0110100100011" => q_unbuf <= my_rom(3363);
      when "0110100100100" => q_unbuf <= my_rom(3364);
      when "0110100100101" => q_unbuf <= my_rom(3365);
      when "0110100100110" => q_unbuf <= my_rom(3366);
      when "0110100100111" => q_unbuf <= my_rom(3367);
      when "0110100101000" => q_unbuf <= my_rom(3368);
      when "0110100101001" => q_unbuf <= my_rom(3369);
      when "0110100101010" => q_unbuf <= my_rom(3370);
      when "0110100101011" => q_unbuf <= my_rom(3371);
      when "0110100101100" => q_unbuf <= my_rom(3372);
      when "0110100101101" => q_unbuf <= my_rom(3373);
      when "0110100101110" => q_unbuf <= my_rom(3374);
      when "0110100101111" => q_unbuf <= my_rom(3375);
      when "0110100110000" => q_unbuf <= my_rom(3376);
      when "0110100110001" => q_unbuf <= my_rom(3377);
      when "0110100110010" => q_unbuf <= my_rom(3378);
      when "0110100110011" => q_unbuf <= my_rom(3379);
      when "0110100110100" => q_unbuf <= my_rom(3380);
      when "0110100110101" => q_unbuf <= my_rom(3381);
      when "0110100110110" => q_unbuf <= my_rom(3382);
      when "0110100110111" => q_unbuf <= my_rom(3383);
      when "0110100111000" => q_unbuf <= my_rom(3384);
      when "0110100111001" => q_unbuf <= my_rom(3385);
      when "0110100111010" => q_unbuf <= my_rom(3386);
      when "0110100111011" => q_unbuf <= my_rom(3387);
      when "0110100111100" => q_unbuf <= my_rom(3388);
      when "0110100111101" => q_unbuf <= my_rom(3389);
      when "0110100111110" => q_unbuf <= my_rom(3390);
      when "0110100111111" => q_unbuf <= my_rom(3391);
      when "0110101000000" => q_unbuf <= my_rom(3392);
      when "0110101000001" => q_unbuf <= my_rom(3393);
      when "0110101000010" => q_unbuf <= my_rom(3394);
      when "0110101000011" => q_unbuf <= my_rom(3395);
      when "0110101000100" => q_unbuf <= my_rom(3396);
      when "0110101000101" => q_unbuf <= my_rom(3397);
      when "0110101000110" => q_unbuf <= my_rom(3398);
      when "0110101000111" => q_unbuf <= my_rom(3399);
      when "0110101001000" => q_unbuf <= my_rom(3400);
      when "0110101001001" => q_unbuf <= my_rom(3401);
      when "0110101001010" => q_unbuf <= my_rom(3402);
      when "0110101001011" => q_unbuf <= my_rom(3403);
      when "0110101001100" => q_unbuf <= my_rom(3404);
      when "0110101001101" => q_unbuf <= my_rom(3405);
      when "0110101001110" => q_unbuf <= my_rom(3406);
      when "0110101001111" => q_unbuf <= my_rom(3407);
      when "0110101010000" => q_unbuf <= my_rom(3408);
      when "0110101010001" => q_unbuf <= my_rom(3409);
      when "0110101010010" => q_unbuf <= my_rom(3410);
      when "0110101010011" => q_unbuf <= my_rom(3411);
      when "0110101010100" => q_unbuf <= my_rom(3412);
      when "0110101010101" => q_unbuf <= my_rom(3413);
      when "0110101010110" => q_unbuf <= my_rom(3414);
      when "0110101010111" => q_unbuf <= my_rom(3415);
      when "0110101011000" => q_unbuf <= my_rom(3416);
      when "0110101011001" => q_unbuf <= my_rom(3417);
      when "0110101011010" => q_unbuf <= my_rom(3418);
      when "0110101011011" => q_unbuf <= my_rom(3419);
      when "0110101011100" => q_unbuf <= my_rom(3420);
      when "0110101011101" => q_unbuf <= my_rom(3421);
      when "0110101011110" => q_unbuf <= my_rom(3422);
      when "0110101011111" => q_unbuf <= my_rom(3423);
      when "0110101100000" => q_unbuf <= my_rom(3424);
      when "0110101100001" => q_unbuf <= my_rom(3425);
      when "0110101100010" => q_unbuf <= my_rom(3426);
      when "0110101100011" => q_unbuf <= my_rom(3427);
      when "0110101100100" => q_unbuf <= my_rom(3428);
      when "0110101100101" => q_unbuf <= my_rom(3429);
      when "0110101100110" => q_unbuf <= my_rom(3430);
      when "0110101100111" => q_unbuf <= my_rom(3431);
      when "0110101101000" => q_unbuf <= my_rom(3432);
      when "0110101101001" => q_unbuf <= my_rom(3433);
      when "0110101101010" => q_unbuf <= my_rom(3434);
      when "0110101101011" => q_unbuf <= my_rom(3435);
      when "0110101101100" => q_unbuf <= my_rom(3436);
      when "0110101101101" => q_unbuf <= my_rom(3437);
      when "0110101101110" => q_unbuf <= my_rom(3438);
      when "0110101101111" => q_unbuf <= my_rom(3439);
      when "0110101110000" => q_unbuf <= my_rom(3440);
      when "0110101110001" => q_unbuf <= my_rom(3441);
      when "0110101110010" => q_unbuf <= my_rom(3442);
      when "0110101110011" => q_unbuf <= my_rom(3443);
      when "0110101110100" => q_unbuf <= my_rom(3444);
      when "0110101110101" => q_unbuf <= my_rom(3445);
      when "0110101110110" => q_unbuf <= my_rom(3446);
      when "0110101110111" => q_unbuf <= my_rom(3447);
      when "0110101111000" => q_unbuf <= my_rom(3448);
      when "0110101111001" => q_unbuf <= my_rom(3449);
      when "0110101111010" => q_unbuf <= my_rom(3450);
      when "0110101111011" => q_unbuf <= my_rom(3451);
      when "0110101111100" => q_unbuf <= my_rom(3452);
      when "0110101111101" => q_unbuf <= my_rom(3453);
      when "0110101111110" => q_unbuf <= my_rom(3454);
      when "0110101111111" => q_unbuf <= my_rom(3455);
      when "0110110000000" => q_unbuf <= my_rom(3456);
      when "0110110000001" => q_unbuf <= my_rom(3457);
      when "0110110000010" => q_unbuf <= my_rom(3458);
      when "0110110000011" => q_unbuf <= my_rom(3459);
      when "0110110000100" => q_unbuf <= my_rom(3460);
      when "0110110000101" => q_unbuf <= my_rom(3461);
      when "0110110000110" => q_unbuf <= my_rom(3462);
      when "0110110000111" => q_unbuf <= my_rom(3463);
      when "0110110001000" => q_unbuf <= my_rom(3464);
      when "0110110001001" => q_unbuf <= my_rom(3465);
      when "0110110001010" => q_unbuf <= my_rom(3466);
      when "0110110001011" => q_unbuf <= my_rom(3467);
      when "0110110001100" => q_unbuf <= my_rom(3468);
      when "0110110001101" => q_unbuf <= my_rom(3469);
      when "0110110001110" => q_unbuf <= my_rom(3470);
      when "0110110001111" => q_unbuf <= my_rom(3471);
      when "0110110010000" => q_unbuf <= my_rom(3472);
      when "0110110010001" => q_unbuf <= my_rom(3473);
      when "0110110010010" => q_unbuf <= my_rom(3474);
      when "0110110010011" => q_unbuf <= my_rom(3475);
      when "0110110010100" => q_unbuf <= my_rom(3476);
      when "0110110010101" => q_unbuf <= my_rom(3477);
      when "0110110010110" => q_unbuf <= my_rom(3478);
      when "0110110010111" => q_unbuf <= my_rom(3479);
      when "0110110011000" => q_unbuf <= my_rom(3480);
      when "0110110011001" => q_unbuf <= my_rom(3481);
      when "0110110011010" => q_unbuf <= my_rom(3482);
      when "0110110011011" => q_unbuf <= my_rom(3483);
      when "0110110011100" => q_unbuf <= my_rom(3484);
      when "0110110011101" => q_unbuf <= my_rom(3485);
      when "0110110011110" => q_unbuf <= my_rom(3486);
      when "0110110011111" => q_unbuf <= my_rom(3487);
      when "0110110100000" => q_unbuf <= my_rom(3488);
      when "0110110100001" => q_unbuf <= my_rom(3489);
      when "0110110100010" => q_unbuf <= my_rom(3490);
      when "0110110100011" => q_unbuf <= my_rom(3491);
      when "0110110100100" => q_unbuf <= my_rom(3492);
      when "0110110100101" => q_unbuf <= my_rom(3493);
      when "0110110100110" => q_unbuf <= my_rom(3494);
      when "0110110100111" => q_unbuf <= my_rom(3495);
      when "0110110101000" => q_unbuf <= my_rom(3496);
      when "0110110101001" => q_unbuf <= my_rom(3497);
      when "0110110101010" => q_unbuf <= my_rom(3498);
      when "0110110101011" => q_unbuf <= my_rom(3499);
      when "0110110101100" => q_unbuf <= my_rom(3500);
      when "0110110101101" => q_unbuf <= my_rom(3501);
      when "0110110101110" => q_unbuf <= my_rom(3502);
      when "0110110101111" => q_unbuf <= my_rom(3503);
      when "0110110110000" => q_unbuf <= my_rom(3504);
      when "0110110110001" => q_unbuf <= my_rom(3505);
      when "0110110110010" => q_unbuf <= my_rom(3506);
      when "0110110110011" => q_unbuf <= my_rom(3507);
      when "0110110110100" => q_unbuf <= my_rom(3508);
      when "0110110110101" => q_unbuf <= my_rom(3509);
      when "0110110110110" => q_unbuf <= my_rom(3510);
      when "0110110110111" => q_unbuf <= my_rom(3511);
      when "0110110111000" => q_unbuf <= my_rom(3512);
      when "0110110111001" => q_unbuf <= my_rom(3513);
      when "0110110111010" => q_unbuf <= my_rom(3514);
      when "0110110111011" => q_unbuf <= my_rom(3515);
      when "0110110111100" => q_unbuf <= my_rom(3516);
      when "0110110111101" => q_unbuf <= my_rom(3517);
      when "0110110111110" => q_unbuf <= my_rom(3518);
      when "0110110111111" => q_unbuf <= my_rom(3519);
      when "0110111000000" => q_unbuf <= my_rom(3520);
      when "0110111000001" => q_unbuf <= my_rom(3521);
      when "0110111000010" => q_unbuf <= my_rom(3522);
      when "0110111000011" => q_unbuf <= my_rom(3523);
      when "0110111000100" => q_unbuf <= my_rom(3524);
      when "0110111000101" => q_unbuf <= my_rom(3525);
      when "0110111000110" => q_unbuf <= my_rom(3526);
      when "0110111000111" => q_unbuf <= my_rom(3527);
      when "0110111001000" => q_unbuf <= my_rom(3528);
      when "0110111001001" => q_unbuf <= my_rom(3529);
      when "0110111001010" => q_unbuf <= my_rom(3530);
      when "0110111001011" => q_unbuf <= my_rom(3531);
      when "0110111001100" => q_unbuf <= my_rom(3532);
      when "0110111001101" => q_unbuf <= my_rom(3533);
      when "0110111001110" => q_unbuf <= my_rom(3534);
      when "0110111001111" => q_unbuf <= my_rom(3535);
      when "0110111010000" => q_unbuf <= my_rom(3536);
      when "0110111010001" => q_unbuf <= my_rom(3537);
      when "0110111010010" => q_unbuf <= my_rom(3538);
      when "0110111010011" => q_unbuf <= my_rom(3539);
      when "0110111010100" => q_unbuf <= my_rom(3540);
      when "0110111010101" => q_unbuf <= my_rom(3541);
      when "0110111010110" => q_unbuf <= my_rom(3542);
      when "0110111010111" => q_unbuf <= my_rom(3543);
      when "0110111011000" => q_unbuf <= my_rom(3544);
      when "0110111011001" => q_unbuf <= my_rom(3545);
      when "0110111011010" => q_unbuf <= my_rom(3546);
      when "0110111011011" => q_unbuf <= my_rom(3547);
      when "0110111011100" => q_unbuf <= my_rom(3548);
      when "0110111011101" => q_unbuf <= my_rom(3549);
      when "0110111011110" => q_unbuf <= my_rom(3550);
      when "0110111011111" => q_unbuf <= my_rom(3551);
      when "0110111100000" => q_unbuf <= my_rom(3552);
      when "0110111100001" => q_unbuf <= my_rom(3553);
      when "0110111100010" => q_unbuf <= my_rom(3554);
      when "0110111100011" => q_unbuf <= my_rom(3555);
      when "0110111100100" => q_unbuf <= my_rom(3556);
      when "0110111100101" => q_unbuf <= my_rom(3557);
      when "0110111100110" => q_unbuf <= my_rom(3558);
      when "0110111100111" => q_unbuf <= my_rom(3559);
      when "0110111101000" => q_unbuf <= my_rom(3560);
      when "0110111101001" => q_unbuf <= my_rom(3561);
      when "0110111101010" => q_unbuf <= my_rom(3562);
      when "0110111101011" => q_unbuf <= my_rom(3563);
      when "0110111101100" => q_unbuf <= my_rom(3564);
      when "0110111101101" => q_unbuf <= my_rom(3565);
      when "0110111101110" => q_unbuf <= my_rom(3566);
      when "0110111101111" => q_unbuf <= my_rom(3567);
      when "0110111110000" => q_unbuf <= my_rom(3568);
      when "0110111110001" => q_unbuf <= my_rom(3569);
      when "0110111110010" => q_unbuf <= my_rom(3570);
      when "0110111110011" => q_unbuf <= my_rom(3571);
      when "0110111110100" => q_unbuf <= my_rom(3572);
      when "0110111110101" => q_unbuf <= my_rom(3573);
      when "0110111110110" => q_unbuf <= my_rom(3574);
      when "0110111110111" => q_unbuf <= my_rom(3575);
      when "0110111111000" => q_unbuf <= my_rom(3576);
      when "0110111111001" => q_unbuf <= my_rom(3577);
      when "0110111111010" => q_unbuf <= my_rom(3578);
      when "0110111111011" => q_unbuf <= my_rom(3579);
      when "0110111111100" => q_unbuf <= my_rom(3580);
      when "0110111111101" => q_unbuf <= my_rom(3581);
      when "0110111111110" => q_unbuf <= my_rom(3582);
      when "0110111111111" => q_unbuf <= my_rom(3583);
      when "0111000000000" => q_unbuf <= my_rom(3584);
      when "0111000000001" => q_unbuf <= my_rom(3585);
      when "0111000000010" => q_unbuf <= my_rom(3586);
      when "0111000000011" => q_unbuf <= my_rom(3587);
      when "0111000000100" => q_unbuf <= my_rom(3588);
      when "0111000000101" => q_unbuf <= my_rom(3589);
      when "0111000000110" => q_unbuf <= my_rom(3590);
      when "0111000000111" => q_unbuf <= my_rom(3591);
      when "0111000001000" => q_unbuf <= my_rom(3592);
      when "0111000001001" => q_unbuf <= my_rom(3593);
      when "0111000001010" => q_unbuf <= my_rom(3594);
      when "0111000001011" => q_unbuf <= my_rom(3595);
      when "0111000001100" => q_unbuf <= my_rom(3596);
      when "0111000001101" => q_unbuf <= my_rom(3597);
      when "0111000001110" => q_unbuf <= my_rom(3598);
      when "0111000001111" => q_unbuf <= my_rom(3599);
      when "0111000010000" => q_unbuf <= my_rom(3600);
      when "0111000010001" => q_unbuf <= my_rom(3601);
      when "0111000010010" => q_unbuf <= my_rom(3602);
      when "0111000010011" => q_unbuf <= my_rom(3603);
      when "0111000010100" => q_unbuf <= my_rom(3604);
      when "0111000010101" => q_unbuf <= my_rom(3605);
      when "0111000010110" => q_unbuf <= my_rom(3606);
      when "0111000010111" => q_unbuf <= my_rom(3607);
      when "0111000011000" => q_unbuf <= my_rom(3608);
      when "0111000011001" => q_unbuf <= my_rom(3609);
      when "0111000011010" => q_unbuf <= my_rom(3610);
      when "0111000011011" => q_unbuf <= my_rom(3611);
      when "0111000011100" => q_unbuf <= my_rom(3612);
      when "0111000011101" => q_unbuf <= my_rom(3613);
      when "0111000011110" => q_unbuf <= my_rom(3614);
      when "0111000011111" => q_unbuf <= my_rom(3615);
      when "0111000100000" => q_unbuf <= my_rom(3616);
      when "0111000100001" => q_unbuf <= my_rom(3617);
      when "0111000100010" => q_unbuf <= my_rom(3618);
      when "0111000100011" => q_unbuf <= my_rom(3619);
      when "0111000100100" => q_unbuf <= my_rom(3620);
      when "0111000100101" => q_unbuf <= my_rom(3621);
      when "0111000100110" => q_unbuf <= my_rom(3622);
      when "0111000100111" => q_unbuf <= my_rom(3623);
      when "0111000101000" => q_unbuf <= my_rom(3624);
      when "0111000101001" => q_unbuf <= my_rom(3625);
      when "0111000101010" => q_unbuf <= my_rom(3626);
      when "0111000101011" => q_unbuf <= my_rom(3627);
      when "0111000101100" => q_unbuf <= my_rom(3628);
      when "0111000101101" => q_unbuf <= my_rom(3629);
      when "0111000101110" => q_unbuf <= my_rom(3630);
      when "0111000101111" => q_unbuf <= my_rom(3631);
      when "0111000110000" => q_unbuf <= my_rom(3632);
      when "0111000110001" => q_unbuf <= my_rom(3633);
      when "0111000110010" => q_unbuf <= my_rom(3634);
      when "0111000110011" => q_unbuf <= my_rom(3635);
      when "0111000110100" => q_unbuf <= my_rom(3636);
      when "0111000110101" => q_unbuf <= my_rom(3637);
      when "0111000110110" => q_unbuf <= my_rom(3638);
      when "0111000110111" => q_unbuf <= my_rom(3639);
      when "0111000111000" => q_unbuf <= my_rom(3640);
      when "0111000111001" => q_unbuf <= my_rom(3641);
      when "0111000111010" => q_unbuf <= my_rom(3642);
      when "0111000111011" => q_unbuf <= my_rom(3643);
      when "0111000111100" => q_unbuf <= my_rom(3644);
      when "0111000111101" => q_unbuf <= my_rom(3645);
      when "0111000111110" => q_unbuf <= my_rom(3646);
      when "0111000111111" => q_unbuf <= my_rom(3647);
      when "0111001000000" => q_unbuf <= my_rom(3648);
      when "0111001000001" => q_unbuf <= my_rom(3649);
      when "0111001000010" => q_unbuf <= my_rom(3650);
      when "0111001000011" => q_unbuf <= my_rom(3651);
      when "0111001000100" => q_unbuf <= my_rom(3652);
      when "0111001000101" => q_unbuf <= my_rom(3653);
      when "0111001000110" => q_unbuf <= my_rom(3654);
      when "0111001000111" => q_unbuf <= my_rom(3655);
      when "0111001001000" => q_unbuf <= my_rom(3656);
      when "0111001001001" => q_unbuf <= my_rom(3657);
      when "0111001001010" => q_unbuf <= my_rom(3658);
      when "0111001001011" => q_unbuf <= my_rom(3659);
      when "0111001001100" => q_unbuf <= my_rom(3660);
      when "0111001001101" => q_unbuf <= my_rom(3661);
      when "0111001001110" => q_unbuf <= my_rom(3662);
      when "0111001001111" => q_unbuf <= my_rom(3663);
      when "0111001010000" => q_unbuf <= my_rom(3664);
      when "0111001010001" => q_unbuf <= my_rom(3665);
      when "0111001010010" => q_unbuf <= my_rom(3666);
      when "0111001010011" => q_unbuf <= my_rom(3667);
      when "0111001010100" => q_unbuf <= my_rom(3668);
      when "0111001010101" => q_unbuf <= my_rom(3669);
      when "0111001010110" => q_unbuf <= my_rom(3670);
      when "0111001010111" => q_unbuf <= my_rom(3671);
      when "0111001011000" => q_unbuf <= my_rom(3672);
      when "0111001011001" => q_unbuf <= my_rom(3673);
      when "0111001011010" => q_unbuf <= my_rom(3674);
      when "0111001011011" => q_unbuf <= my_rom(3675);
      when "0111001011100" => q_unbuf <= my_rom(3676);
      when "0111001011101" => q_unbuf <= my_rom(3677);
      when "0111001011110" => q_unbuf <= my_rom(3678);
      when "0111001011111" => q_unbuf <= my_rom(3679);
      when "0111001100000" => q_unbuf <= my_rom(3680);
      when "0111001100001" => q_unbuf <= my_rom(3681);
      when "0111001100010" => q_unbuf <= my_rom(3682);
      when "0111001100011" => q_unbuf <= my_rom(3683);
      when "0111001100100" => q_unbuf <= my_rom(3684);
      when "0111001100101" => q_unbuf <= my_rom(3685);
      when "0111001100110" => q_unbuf <= my_rom(3686);
      when "0111001100111" => q_unbuf <= my_rom(3687);
      when "0111001101000" => q_unbuf <= my_rom(3688);
      when "0111001101001" => q_unbuf <= my_rom(3689);
      when "0111001101010" => q_unbuf <= my_rom(3690);
      when "0111001101011" => q_unbuf <= my_rom(3691);
      when "0111001101100" => q_unbuf <= my_rom(3692);
      when "0111001101101" => q_unbuf <= my_rom(3693);
      when "0111001101110" => q_unbuf <= my_rom(3694);
      when "0111001101111" => q_unbuf <= my_rom(3695);
      when "0111001110000" => q_unbuf <= my_rom(3696);
      when "0111001110001" => q_unbuf <= my_rom(3697);
      when "0111001110010" => q_unbuf <= my_rom(3698);
      when "0111001110011" => q_unbuf <= my_rom(3699);
      when "0111001110100" => q_unbuf <= my_rom(3700);
      when "0111001110101" => q_unbuf <= my_rom(3701);
      when "0111001110110" => q_unbuf <= my_rom(3702);
      when "0111001110111" => q_unbuf <= my_rom(3703);
      when "0111001111000" => q_unbuf <= my_rom(3704);
      when "0111001111001" => q_unbuf <= my_rom(3705);
      when "0111001111010" => q_unbuf <= my_rom(3706);
      when "0111001111011" => q_unbuf <= my_rom(3707);
      when "0111001111100" => q_unbuf <= my_rom(3708);
      when "0111001111101" => q_unbuf <= my_rom(3709);
      when "0111001111110" => q_unbuf <= my_rom(3710);
      when "0111001111111" => q_unbuf <= my_rom(3711);
      when "0111010000000" => q_unbuf <= my_rom(3712);
      when "0111010000001" => q_unbuf <= my_rom(3713);
      when "0111010000010" => q_unbuf <= my_rom(3714);
      when "0111010000011" => q_unbuf <= my_rom(3715);
      when "0111010000100" => q_unbuf <= my_rom(3716);
      when "0111010000101" => q_unbuf <= my_rom(3717);
      when "0111010000110" => q_unbuf <= my_rom(3718);
      when "0111010000111" => q_unbuf <= my_rom(3719);
      when "0111010001000" => q_unbuf <= my_rom(3720);
      when "0111010001001" => q_unbuf <= my_rom(3721);
      when "0111010001010" => q_unbuf <= my_rom(3722);
      when "0111010001011" => q_unbuf <= my_rom(3723);
      when "0111010001100" => q_unbuf <= my_rom(3724);
      when "0111010001101" => q_unbuf <= my_rom(3725);
      when "0111010001110" => q_unbuf <= my_rom(3726);
      when "0111010001111" => q_unbuf <= my_rom(3727);
      when "0111010010000" => q_unbuf <= my_rom(3728);
      when "0111010010001" => q_unbuf <= my_rom(3729);
      when "0111010010010" => q_unbuf <= my_rom(3730);
      when "0111010010011" => q_unbuf <= my_rom(3731);
      when "0111010010100" => q_unbuf <= my_rom(3732);
      when "0111010010101" => q_unbuf <= my_rom(3733);
      when "0111010010110" => q_unbuf <= my_rom(3734);
      when "0111010010111" => q_unbuf <= my_rom(3735);
      when "0111010011000" => q_unbuf <= my_rom(3736);
      when "0111010011001" => q_unbuf <= my_rom(3737);
      when "0111010011010" => q_unbuf <= my_rom(3738);
      when "0111010011011" => q_unbuf <= my_rom(3739);
      when "0111010011100" => q_unbuf <= my_rom(3740);
      when "0111010011101" => q_unbuf <= my_rom(3741);
      when "0111010011110" => q_unbuf <= my_rom(3742);
      when "0111010011111" => q_unbuf <= my_rom(3743);
      when "0111010100000" => q_unbuf <= my_rom(3744);
      when "0111010100001" => q_unbuf <= my_rom(3745);
      when "0111010100010" => q_unbuf <= my_rom(3746);
      when "0111010100011" => q_unbuf <= my_rom(3747);
      when "0111010100100" => q_unbuf <= my_rom(3748);
      when "0111010100101" => q_unbuf <= my_rom(3749);
      when "0111010100110" => q_unbuf <= my_rom(3750);
      when "0111010100111" => q_unbuf <= my_rom(3751);
      when "0111010101000" => q_unbuf <= my_rom(3752);
      when "0111010101001" => q_unbuf <= my_rom(3753);
      when "0111010101010" => q_unbuf <= my_rom(3754);
      when "0111010101011" => q_unbuf <= my_rom(3755);
      when "0111010101100" => q_unbuf <= my_rom(3756);
      when "0111010101101" => q_unbuf <= my_rom(3757);
      when "0111010101110" => q_unbuf <= my_rom(3758);
      when "0111010101111" => q_unbuf <= my_rom(3759);
      when "0111010110000" => q_unbuf <= my_rom(3760);
      when "0111010110001" => q_unbuf <= my_rom(3761);
      when "0111010110010" => q_unbuf <= my_rom(3762);
      when "0111010110011" => q_unbuf <= my_rom(3763);
      when "0111010110100" => q_unbuf <= my_rom(3764);
      when "0111010110101" => q_unbuf <= my_rom(3765);
      when "0111010110110" => q_unbuf <= my_rom(3766);
      when "0111010110111" => q_unbuf <= my_rom(3767);
      when "0111010111000" => q_unbuf <= my_rom(3768);
      when "0111010111001" => q_unbuf <= my_rom(3769);
      when "0111010111010" => q_unbuf <= my_rom(3770);
      when "0111010111011" => q_unbuf <= my_rom(3771);
      when "0111010111100" => q_unbuf <= my_rom(3772);
      when "0111010111101" => q_unbuf <= my_rom(3773);
      when "0111010111110" => q_unbuf <= my_rom(3774);
      when "0111010111111" => q_unbuf <= my_rom(3775);
      when "0111011000000" => q_unbuf <= my_rom(3776);
      when "0111011000001" => q_unbuf <= my_rom(3777);
      when "0111011000010" => q_unbuf <= my_rom(3778);
      when "0111011000011" => q_unbuf <= my_rom(3779);
      when "0111011000100" => q_unbuf <= my_rom(3780);
      when "0111011000101" => q_unbuf <= my_rom(3781);
      when "0111011000110" => q_unbuf <= my_rom(3782);
      when "0111011000111" => q_unbuf <= my_rom(3783);
      when "0111011001000" => q_unbuf <= my_rom(3784);
      when "0111011001001" => q_unbuf <= my_rom(3785);
      when "0111011001010" => q_unbuf <= my_rom(3786);
      when "0111011001011" => q_unbuf <= my_rom(3787);
      when "0111011001100" => q_unbuf <= my_rom(3788);
      when "0111011001101" => q_unbuf <= my_rom(3789);
      when "0111011001110" => q_unbuf <= my_rom(3790);
      when "0111011001111" => q_unbuf <= my_rom(3791);
      when "0111011010000" => q_unbuf <= my_rom(3792);
      when "0111011010001" => q_unbuf <= my_rom(3793);
      when "0111011010010" => q_unbuf <= my_rom(3794);
      when "0111011010011" => q_unbuf <= my_rom(3795);
      when "0111011010100" => q_unbuf <= my_rom(3796);
      when "0111011010101" => q_unbuf <= my_rom(3797);
      when "0111011010110" => q_unbuf <= my_rom(3798);
      when "0111011010111" => q_unbuf <= my_rom(3799);
      when "0111011011000" => q_unbuf <= my_rom(3800);
      when "0111011011001" => q_unbuf <= my_rom(3801);
      when "0111011011010" => q_unbuf <= my_rom(3802);
      when "0111011011011" => q_unbuf <= my_rom(3803);
      when "0111011011100" => q_unbuf <= my_rom(3804);
      when "0111011011101" => q_unbuf <= my_rom(3805);
      when "0111011011110" => q_unbuf <= my_rom(3806);
      when "0111011011111" => q_unbuf <= my_rom(3807);
      when "0111011100000" => q_unbuf <= my_rom(3808);
      when "0111011100001" => q_unbuf <= my_rom(3809);
      when "0111011100010" => q_unbuf <= my_rom(3810);
      when "0111011100011" => q_unbuf <= my_rom(3811);
      when "0111011100100" => q_unbuf <= my_rom(3812);
      when "0111011100101" => q_unbuf <= my_rom(3813);
      when "0111011100110" => q_unbuf <= my_rom(3814);
      when "0111011100111" => q_unbuf <= my_rom(3815);
      when "0111011101000" => q_unbuf <= my_rom(3816);
      when "0111011101001" => q_unbuf <= my_rom(3817);
      when "0111011101010" => q_unbuf <= my_rom(3818);
      when "0111011101011" => q_unbuf <= my_rom(3819);
      when "0111011101100" => q_unbuf <= my_rom(3820);
      when "0111011101101" => q_unbuf <= my_rom(3821);
      when "0111011101110" => q_unbuf <= my_rom(3822);
      when "0111011101111" => q_unbuf <= my_rom(3823);
      when "0111011110000" => q_unbuf <= my_rom(3824);
      when "0111011110001" => q_unbuf <= my_rom(3825);
      when "0111011110010" => q_unbuf <= my_rom(3826);
      when "0111011110011" => q_unbuf <= my_rom(3827);
      when "0111011110100" => q_unbuf <= my_rom(3828);
      when "0111011110101" => q_unbuf <= my_rom(3829);
      when "0111011110110" => q_unbuf <= my_rom(3830);
      when "0111011110111" => q_unbuf <= my_rom(3831);
      when "0111011111000" => q_unbuf <= my_rom(3832);
      when "0111011111001" => q_unbuf <= my_rom(3833);
      when "0111011111010" => q_unbuf <= my_rom(3834);
      when "0111011111011" => q_unbuf <= my_rom(3835);
      when "0111011111100" => q_unbuf <= my_rom(3836);
      when "0111011111101" => q_unbuf <= my_rom(3837);
      when "0111011111110" => q_unbuf <= my_rom(3838);
      when "0111011111111" => q_unbuf <= my_rom(3839);
      when "0111100000000" => q_unbuf <= my_rom(3840);
      when "0111100000001" => q_unbuf <= my_rom(3841);
      when "0111100000010" => q_unbuf <= my_rom(3842);
      when "0111100000011" => q_unbuf <= my_rom(3843);
      when "0111100000100" => q_unbuf <= my_rom(3844);
      when "0111100000101" => q_unbuf <= my_rom(3845);
      when "0111100000110" => q_unbuf <= my_rom(3846);
      when "0111100000111" => q_unbuf <= my_rom(3847);
      when "0111100001000" => q_unbuf <= my_rom(3848);
      when "0111100001001" => q_unbuf <= my_rom(3849);
      when "0111100001010" => q_unbuf <= my_rom(3850);
      when "0111100001011" => q_unbuf <= my_rom(3851);
      when "0111100001100" => q_unbuf <= my_rom(3852);
      when "0111100001101" => q_unbuf <= my_rom(3853);
      when "0111100001110" => q_unbuf <= my_rom(3854);
      when "0111100001111" => q_unbuf <= my_rom(3855);
      when "0111100010000" => q_unbuf <= my_rom(3856);
      when "0111100010001" => q_unbuf <= my_rom(3857);
      when "0111100010010" => q_unbuf <= my_rom(3858);
      when "0111100010011" => q_unbuf <= my_rom(3859);
      when "0111100010100" => q_unbuf <= my_rom(3860);
      when "0111100010101" => q_unbuf <= my_rom(3861);
      when "0111100010110" => q_unbuf <= my_rom(3862);
      when "0111100010111" => q_unbuf <= my_rom(3863);
      when "0111100011000" => q_unbuf <= my_rom(3864);
      when "0111100011001" => q_unbuf <= my_rom(3865);
      when "0111100011010" => q_unbuf <= my_rom(3866);
      when "0111100011011" => q_unbuf <= my_rom(3867);
      when "0111100011100" => q_unbuf <= my_rom(3868);
      when "0111100011101" => q_unbuf <= my_rom(3869);
      when "0111100011110" => q_unbuf <= my_rom(3870);
      when "0111100011111" => q_unbuf <= my_rom(3871);
      when "0111100100000" => q_unbuf <= my_rom(3872);
      when "0111100100001" => q_unbuf <= my_rom(3873);
      when "0111100100010" => q_unbuf <= my_rom(3874);
      when "0111100100011" => q_unbuf <= my_rom(3875);
      when "0111100100100" => q_unbuf <= my_rom(3876);
      when "0111100100101" => q_unbuf <= my_rom(3877);
      when "0111100100110" => q_unbuf <= my_rom(3878);
      when "0111100100111" => q_unbuf <= my_rom(3879);
      when "0111100101000" => q_unbuf <= my_rom(3880);
      when "0111100101001" => q_unbuf <= my_rom(3881);
      when "0111100101010" => q_unbuf <= my_rom(3882);
      when "0111100101011" => q_unbuf <= my_rom(3883);
      when "0111100101100" => q_unbuf <= my_rom(3884);
      when "0111100101101" => q_unbuf <= my_rom(3885);
      when "0111100101110" => q_unbuf <= my_rom(3886);
      when "0111100101111" => q_unbuf <= my_rom(3887);
      when "0111100110000" => q_unbuf <= my_rom(3888);
      when "0111100110001" => q_unbuf <= my_rom(3889);
      when "0111100110010" => q_unbuf <= my_rom(3890);
      when "0111100110011" => q_unbuf <= my_rom(3891);
      when "0111100110100" => q_unbuf <= my_rom(3892);
      when "0111100110101" => q_unbuf <= my_rom(3893);
      when "0111100110110" => q_unbuf <= my_rom(3894);
      when "0111100110111" => q_unbuf <= my_rom(3895);
      when "0111100111000" => q_unbuf <= my_rom(3896);
      when "0111100111001" => q_unbuf <= my_rom(3897);
      when "0111100111010" => q_unbuf <= my_rom(3898);
      when "0111100111011" => q_unbuf <= my_rom(3899);
      when "0111100111100" => q_unbuf <= my_rom(3900);
      when "0111100111101" => q_unbuf <= my_rom(3901);
      when "0111100111110" => q_unbuf <= my_rom(3902);
      when "0111100111111" => q_unbuf <= my_rom(3903);
      when "0111101000000" => q_unbuf <= my_rom(3904);
      when "0111101000001" => q_unbuf <= my_rom(3905);
      when "0111101000010" => q_unbuf <= my_rom(3906);
      when "0111101000011" => q_unbuf <= my_rom(3907);
      when "0111101000100" => q_unbuf <= my_rom(3908);
      when "0111101000101" => q_unbuf <= my_rom(3909);
      when "0111101000110" => q_unbuf <= my_rom(3910);
      when "0111101000111" => q_unbuf <= my_rom(3911);
      when "0111101001000" => q_unbuf <= my_rom(3912);
      when "0111101001001" => q_unbuf <= my_rom(3913);
      when "0111101001010" => q_unbuf <= my_rom(3914);
      when "0111101001011" => q_unbuf <= my_rom(3915);
      when "0111101001100" => q_unbuf <= my_rom(3916);
      when "0111101001101" => q_unbuf <= my_rom(3917);
      when "0111101001110" => q_unbuf <= my_rom(3918);
      when "0111101001111" => q_unbuf <= my_rom(3919);
      when "0111101010000" => q_unbuf <= my_rom(3920);
      when "0111101010001" => q_unbuf <= my_rom(3921);
      when "0111101010010" => q_unbuf <= my_rom(3922);
      when "0111101010011" => q_unbuf <= my_rom(3923);
      when "0111101010100" => q_unbuf <= my_rom(3924);
      when "0111101010101" => q_unbuf <= my_rom(3925);
      when "0111101010110" => q_unbuf <= my_rom(3926);
      when "0111101010111" => q_unbuf <= my_rom(3927);
      when "0111101011000" => q_unbuf <= my_rom(3928);
      when "0111101011001" => q_unbuf <= my_rom(3929);
      when "0111101011010" => q_unbuf <= my_rom(3930);
      when "0111101011011" => q_unbuf <= my_rom(3931);
      when "0111101011100" => q_unbuf <= my_rom(3932);
      when "0111101011101" => q_unbuf <= my_rom(3933);
      when "0111101011110" => q_unbuf <= my_rom(3934);
      when "0111101011111" => q_unbuf <= my_rom(3935);
      when "0111101100000" => q_unbuf <= my_rom(3936);
      when "0111101100001" => q_unbuf <= my_rom(3937);
      when "0111101100010" => q_unbuf <= my_rom(3938);
      when "0111101100011" => q_unbuf <= my_rom(3939);
      when "0111101100100" => q_unbuf <= my_rom(3940);
      when "0111101100101" => q_unbuf <= my_rom(3941);
      when "0111101100110" => q_unbuf <= my_rom(3942);
      when "0111101100111" => q_unbuf <= my_rom(3943);
      when "0111101101000" => q_unbuf <= my_rom(3944);
      when "0111101101001" => q_unbuf <= my_rom(3945);
      when "0111101101010" => q_unbuf <= my_rom(3946);
      when "0111101101011" => q_unbuf <= my_rom(3947);
      when "0111101101100" => q_unbuf <= my_rom(3948);
      when "0111101101101" => q_unbuf <= my_rom(3949);
      when "0111101101110" => q_unbuf <= my_rom(3950);
      when "0111101101111" => q_unbuf <= my_rom(3951);
      when "0111101110000" => q_unbuf <= my_rom(3952);
      when "0111101110001" => q_unbuf <= my_rom(3953);
      when "0111101110010" => q_unbuf <= my_rom(3954);
      when "0111101110011" => q_unbuf <= my_rom(3955);
      when "0111101110100" => q_unbuf <= my_rom(3956);
      when "0111101110101" => q_unbuf <= my_rom(3957);
      when "0111101110110" => q_unbuf <= my_rom(3958);
      when "0111101110111" => q_unbuf <= my_rom(3959);
      when "0111101111000" => q_unbuf <= my_rom(3960);
      when "0111101111001" => q_unbuf <= my_rom(3961);
      when "0111101111010" => q_unbuf <= my_rom(3962);
      when "0111101111011" => q_unbuf <= my_rom(3963);
      when "0111101111100" => q_unbuf <= my_rom(3964);
      when "0111101111101" => q_unbuf <= my_rom(3965);
      when "0111101111110" => q_unbuf <= my_rom(3966);
      when "0111101111111" => q_unbuf <= my_rom(3967);
      when "0111110000000" => q_unbuf <= my_rom(3968);
      when "0111110000001" => q_unbuf <= my_rom(3969);
      when "0111110000010" => q_unbuf <= my_rom(3970);
      when "0111110000011" => q_unbuf <= my_rom(3971);
      when "0111110000100" => q_unbuf <= my_rom(3972);
      when "0111110000101" => q_unbuf <= my_rom(3973);
      when "0111110000110" => q_unbuf <= my_rom(3974);
      when "0111110000111" => q_unbuf <= my_rom(3975);
      when "0111110001000" => q_unbuf <= my_rom(3976);
      when "0111110001001" => q_unbuf <= my_rom(3977);
      when "0111110001010" => q_unbuf <= my_rom(3978);
      when "0111110001011" => q_unbuf <= my_rom(3979);
      when "0111110001100" => q_unbuf <= my_rom(3980);
      when "0111110001101" => q_unbuf <= my_rom(3981);
      when "0111110001110" => q_unbuf <= my_rom(3982);
      when "0111110001111" => q_unbuf <= my_rom(3983);
      when "0111110010000" => q_unbuf <= my_rom(3984);
      when "0111110010001" => q_unbuf <= my_rom(3985);
      when "0111110010010" => q_unbuf <= my_rom(3986);
      when "0111110010011" => q_unbuf <= my_rom(3987);
      when "0111110010100" => q_unbuf <= my_rom(3988);
      when "0111110010101" => q_unbuf <= my_rom(3989);
      when "0111110010110" => q_unbuf <= my_rom(3990);
      when "0111110010111" => q_unbuf <= my_rom(3991);
      when "0111110011000" => q_unbuf <= my_rom(3992);
      when "0111110011001" => q_unbuf <= my_rom(3993);
      when "0111110011010" => q_unbuf <= my_rom(3994);
      when "0111110011011" => q_unbuf <= my_rom(3995);
      when "0111110011100" => q_unbuf <= my_rom(3996);
      when "0111110011101" => q_unbuf <= my_rom(3997);
      when "0111110011110" => q_unbuf <= my_rom(3998);
      when "0111110011111" => q_unbuf <= my_rom(3999);
      when "0111110100000" => q_unbuf <= my_rom(4000);
      when "0111110100001" => q_unbuf <= my_rom(4001);
      when "0111110100010" => q_unbuf <= my_rom(4002);
      when "0111110100011" => q_unbuf <= my_rom(4003);
      when "0111110100100" => q_unbuf <= my_rom(4004);
      when "0111110100101" => q_unbuf <= my_rom(4005);
      when "0111110100110" => q_unbuf <= my_rom(4006);
      when "0111110100111" => q_unbuf <= my_rom(4007);
      when "0111110101000" => q_unbuf <= my_rom(4008);
      when "0111110101001" => q_unbuf <= my_rom(4009);
      when "0111110101010" => q_unbuf <= my_rom(4010);
      when "0111110101011" => q_unbuf <= my_rom(4011);
      when "0111110101100" => q_unbuf <= my_rom(4012);
      when "0111110101101" => q_unbuf <= my_rom(4013);
      when "0111110101110" => q_unbuf <= my_rom(4014);
      when "0111110101111" => q_unbuf <= my_rom(4015);
      when "0111110110000" => q_unbuf <= my_rom(4016);
      when "0111110110001" => q_unbuf <= my_rom(4017);
      when "0111110110010" => q_unbuf <= my_rom(4018);
      when "0111110110011" => q_unbuf <= my_rom(4019);
      when "0111110110100" => q_unbuf <= my_rom(4020);
      when "0111110110101" => q_unbuf <= my_rom(4021);
      when "0111110110110" => q_unbuf <= my_rom(4022);
      when "0111110110111" => q_unbuf <= my_rom(4023);
      when "0111110111000" => q_unbuf <= my_rom(4024);
      when "0111110111001" => q_unbuf <= my_rom(4025);
      when "0111110111010" => q_unbuf <= my_rom(4026);
      when "0111110111011" => q_unbuf <= my_rom(4027);
      when "0111110111100" => q_unbuf <= my_rom(4028);
      when "0111110111101" => q_unbuf <= my_rom(4029);
      when "0111110111110" => q_unbuf <= my_rom(4030);
      when "0111110111111" => q_unbuf <= my_rom(4031);
      when "0111111000000" => q_unbuf <= my_rom(4032);
      when "0111111000001" => q_unbuf <= my_rom(4033);
      when "0111111000010" => q_unbuf <= my_rom(4034);
      when "0111111000011" => q_unbuf <= my_rom(4035);
      when "0111111000100" => q_unbuf <= my_rom(4036);
      when "0111111000101" => q_unbuf <= my_rom(4037);
      when "0111111000110" => q_unbuf <= my_rom(4038);
      when "0111111000111" => q_unbuf <= my_rom(4039);
      when "0111111001000" => q_unbuf <= my_rom(4040);
      when "0111111001001" => q_unbuf <= my_rom(4041);
      when "0111111001010" => q_unbuf <= my_rom(4042);
      when "0111111001011" => q_unbuf <= my_rom(4043);
      when "0111111001100" => q_unbuf <= my_rom(4044);
      when "0111111001101" => q_unbuf <= my_rom(4045);
      when "0111111001110" => q_unbuf <= my_rom(4046);
      when "0111111001111" => q_unbuf <= my_rom(4047);
      when "0111111010000" => q_unbuf <= my_rom(4048);
      when "0111111010001" => q_unbuf <= my_rom(4049);
      when "0111111010010" => q_unbuf <= my_rom(4050);
      when "0111111010011" => q_unbuf <= my_rom(4051);
      when "0111111010100" => q_unbuf <= my_rom(4052);
      when "0111111010101" => q_unbuf <= my_rom(4053);
      when "0111111010110" => q_unbuf <= my_rom(4054);
      when "0111111010111" => q_unbuf <= my_rom(4055);
      when "0111111011000" => q_unbuf <= my_rom(4056);
      when "0111111011001" => q_unbuf <= my_rom(4057);
      when "0111111011010" => q_unbuf <= my_rom(4058);
      when "0111111011011" => q_unbuf <= my_rom(4059);
      when "0111111011100" => q_unbuf <= my_rom(4060);
      when "0111111011101" => q_unbuf <= my_rom(4061);
      when "0111111011110" => q_unbuf <= my_rom(4062);
      when "0111111011111" => q_unbuf <= my_rom(4063);
      when "0111111100000" => q_unbuf <= my_rom(4064);
      when "0111111100001" => q_unbuf <= my_rom(4065);
      when "0111111100010" => q_unbuf <= my_rom(4066);
      when "0111111100011" => q_unbuf <= my_rom(4067);
      when "0111111100100" => q_unbuf <= my_rom(4068);
      when "0111111100101" => q_unbuf <= my_rom(4069);
      when "0111111100110" => q_unbuf <= my_rom(4070);
      when "0111111100111" => q_unbuf <= my_rom(4071);
      when "0111111101000" => q_unbuf <= my_rom(4072);
      when "0111111101001" => q_unbuf <= my_rom(4073);
      when "0111111101010" => q_unbuf <= my_rom(4074);
      when "0111111101011" => q_unbuf <= my_rom(4075);
      when "0111111101100" => q_unbuf <= my_rom(4076);
      when "0111111101101" => q_unbuf <= my_rom(4077);
      when "0111111101110" => q_unbuf <= my_rom(4078);
      when "0111111101111" => q_unbuf <= my_rom(4079);
      when "0111111110000" => q_unbuf <= my_rom(4080);
      when "0111111110001" => q_unbuf <= my_rom(4081);
      when "0111111110010" => q_unbuf <= my_rom(4082);
      when "0111111110011" => q_unbuf <= my_rom(4083);
      when "0111111110100" => q_unbuf <= my_rom(4084);
      when "0111111110101" => q_unbuf <= my_rom(4085);
      when "0111111110110" => q_unbuf <= my_rom(4086);
      when "0111111110111" => q_unbuf <= my_rom(4087);
      when "0111111111000" => q_unbuf <= my_rom(4088);
      when "0111111111001" => q_unbuf <= my_rom(4089);
      when "0111111111010" => q_unbuf <= my_rom(4090);
      when "0111111111011" => q_unbuf <= my_rom(4091);
      when "0111111111100" => q_unbuf <= my_rom(4092);
      when "0111111111101" => q_unbuf <= my_rom(4093);
      when "0111111111110" => q_unbuf <= my_rom(4094);
      when "0111111111111" => q_unbuf <= my_rom(4095);
      when "1000000000000" => q_unbuf <= my_rom(4096);
      when "1000000000001" => q_unbuf <= my_rom(4097);
      when "1000000000010" => q_unbuf <= my_rom(4098);
      when "1000000000011" => q_unbuf <= my_rom(4099);
      when "1000000000100" => q_unbuf <= my_rom(4100);
      when "1000000000101" => q_unbuf <= my_rom(4101);
      when "1000000000110" => q_unbuf <= my_rom(4102);
      when "1000000000111" => q_unbuf <= my_rom(4103);
      when "1000000001000" => q_unbuf <= my_rom(4104);
      when "1000000001001" => q_unbuf <= my_rom(4105);
      when "1000000001010" => q_unbuf <= my_rom(4106);
      when "1000000001011" => q_unbuf <= my_rom(4107);
      when "1000000001100" => q_unbuf <= my_rom(4108);
      when "1000000001101" => q_unbuf <= my_rom(4109);
      when "1000000001110" => q_unbuf <= my_rom(4110);
      when "1000000001111" => q_unbuf <= my_rom(4111);
      when "1000000010000" => q_unbuf <= my_rom(4112);
      when "1000000010001" => q_unbuf <= my_rom(4113);
      when "1000000010010" => q_unbuf <= my_rom(4114);
      when "1000000010011" => q_unbuf <= my_rom(4115);
      when "1000000010100" => q_unbuf <= my_rom(4116);
      when "1000000010101" => q_unbuf <= my_rom(4117);
      when "1000000010110" => q_unbuf <= my_rom(4118);
      when "1000000010111" => q_unbuf <= my_rom(4119);
      when "1000000011000" => q_unbuf <= my_rom(4120);
      when "1000000011001" => q_unbuf <= my_rom(4121);
      when "1000000011010" => q_unbuf <= my_rom(4122);
      when "1000000011011" => q_unbuf <= my_rom(4123);
      when "1000000011100" => q_unbuf <= my_rom(4124);
      when "1000000011101" => q_unbuf <= my_rom(4125);
      when "1000000011110" => q_unbuf <= my_rom(4126);
      when "1000000011111" => q_unbuf <= my_rom(4127);
      when "1000000100000" => q_unbuf <= my_rom(4128);
      when "1000000100001" => q_unbuf <= my_rom(4129);
      when "1000000100010" => q_unbuf <= my_rom(4130);
      when "1000000100011" => q_unbuf <= my_rom(4131);
      when "1000000100100" => q_unbuf <= my_rom(4132);
      when "1000000100101" => q_unbuf <= my_rom(4133);
      when "1000000100110" => q_unbuf <= my_rom(4134);
      when "1000000100111" => q_unbuf <= my_rom(4135);
      when "1000000101000" => q_unbuf <= my_rom(4136);
      when "1000000101001" => q_unbuf <= my_rom(4137);
      when "1000000101010" => q_unbuf <= my_rom(4138);
      when "1000000101011" => q_unbuf <= my_rom(4139);
      when "1000000101100" => q_unbuf <= my_rom(4140);
      when "1000000101101" => q_unbuf <= my_rom(4141);
      when "1000000101110" => q_unbuf <= my_rom(4142);
      when "1000000101111" => q_unbuf <= my_rom(4143);
      when "1000000110000" => q_unbuf <= my_rom(4144);
      when "1000000110001" => q_unbuf <= my_rom(4145);
      when "1000000110010" => q_unbuf <= my_rom(4146);
      when "1000000110011" => q_unbuf <= my_rom(4147);
      when "1000000110100" => q_unbuf <= my_rom(4148);
      when "1000000110101" => q_unbuf <= my_rom(4149);
      when "1000000110110" => q_unbuf <= my_rom(4150);
      when "1000000110111" => q_unbuf <= my_rom(4151);
      when "1000000111000" => q_unbuf <= my_rom(4152);
      when "1000000111001" => q_unbuf <= my_rom(4153);
      when "1000000111010" => q_unbuf <= my_rom(4154);
      when "1000000111011" => q_unbuf <= my_rom(4155);
      when "1000000111100" => q_unbuf <= my_rom(4156);
      when "1000000111101" => q_unbuf <= my_rom(4157);
      when "1000000111110" => q_unbuf <= my_rom(4158);
      when "1000000111111" => q_unbuf <= my_rom(4159);
      when "1000001000000" => q_unbuf <= my_rom(4160);
      when "1000001000001" => q_unbuf <= my_rom(4161);
      when "1000001000010" => q_unbuf <= my_rom(4162);
      when "1000001000011" => q_unbuf <= my_rom(4163);
      when "1000001000100" => q_unbuf <= my_rom(4164);
      when "1000001000101" => q_unbuf <= my_rom(4165);
      when "1000001000110" => q_unbuf <= my_rom(4166);
      when "1000001000111" => q_unbuf <= my_rom(4167);
      when "1000001001000" => q_unbuf <= my_rom(4168);
      when "1000001001001" => q_unbuf <= my_rom(4169);
      when "1000001001010" => q_unbuf <= my_rom(4170);
      when "1000001001011" => q_unbuf <= my_rom(4171);
      when "1000001001100" => q_unbuf <= my_rom(4172);
      when "1000001001101" => q_unbuf <= my_rom(4173);
      when "1000001001110" => q_unbuf <= my_rom(4174);
      when "1000001001111" => q_unbuf <= my_rom(4175);
      when "1000001010000" => q_unbuf <= my_rom(4176);
      when "1000001010001" => q_unbuf <= my_rom(4177);
      when "1000001010010" => q_unbuf <= my_rom(4178);
      when "1000001010011" => q_unbuf <= my_rom(4179);
      when "1000001010100" => q_unbuf <= my_rom(4180);
      when "1000001010101" => q_unbuf <= my_rom(4181);
      when "1000001010110" => q_unbuf <= my_rom(4182);
      when "1000001010111" => q_unbuf <= my_rom(4183);
      when "1000001011000" => q_unbuf <= my_rom(4184);
      when "1000001011001" => q_unbuf <= my_rom(4185);
      when "1000001011010" => q_unbuf <= my_rom(4186);
      when "1000001011011" => q_unbuf <= my_rom(4187);
      when "1000001011100" => q_unbuf <= my_rom(4188);
      when "1000001011101" => q_unbuf <= my_rom(4189);
      when "1000001011110" => q_unbuf <= my_rom(4190);
      when "1000001011111" => q_unbuf <= my_rom(4191);
      when "1000001100000" => q_unbuf <= my_rom(4192);
      when "1000001100001" => q_unbuf <= my_rom(4193);
      when "1000001100010" => q_unbuf <= my_rom(4194);
      when "1000001100011" => q_unbuf <= my_rom(4195);
      when "1000001100100" => q_unbuf <= my_rom(4196);
      when "1000001100101" => q_unbuf <= my_rom(4197);
      when "1000001100110" => q_unbuf <= my_rom(4198);
      when "1000001100111" => q_unbuf <= my_rom(4199);
      when "1000001101000" => q_unbuf <= my_rom(4200);
      when "1000001101001" => q_unbuf <= my_rom(4201);
      when "1000001101010" => q_unbuf <= my_rom(4202);
      when "1000001101011" => q_unbuf <= my_rom(4203);
      when "1000001101100" => q_unbuf <= my_rom(4204);
      when "1000001101101" => q_unbuf <= my_rom(4205);
      when "1000001101110" => q_unbuf <= my_rom(4206);
      when "1000001101111" => q_unbuf <= my_rom(4207);
      when "1000001110000" => q_unbuf <= my_rom(4208);
      when "1000001110001" => q_unbuf <= my_rom(4209);
      when "1000001110010" => q_unbuf <= my_rom(4210);
      when "1000001110011" => q_unbuf <= my_rom(4211);
      when "1000001110100" => q_unbuf <= my_rom(4212);
      when "1000001110101" => q_unbuf <= my_rom(4213);
      when "1000001110110" => q_unbuf <= my_rom(4214);
      when "1000001110111" => q_unbuf <= my_rom(4215);
      when "1000001111000" => q_unbuf <= my_rom(4216);
      when "1000001111001" => q_unbuf <= my_rom(4217);
      when "1000001111010" => q_unbuf <= my_rom(4218);
      when "1000001111011" => q_unbuf <= my_rom(4219);
      when "1000001111100" => q_unbuf <= my_rom(4220);
      when "1000001111101" => q_unbuf <= my_rom(4221);
      when "1000001111110" => q_unbuf <= my_rom(4222);
      when "1000001111111" => q_unbuf <= my_rom(4223);
      when "1000010000000" => q_unbuf <= my_rom(4224);
      when "1000010000001" => q_unbuf <= my_rom(4225);
      when "1000010000010" => q_unbuf <= my_rom(4226);
      when "1000010000011" => q_unbuf <= my_rom(4227);
      when "1000010000100" => q_unbuf <= my_rom(4228);
      when "1000010000101" => q_unbuf <= my_rom(4229);
      when "1000010000110" => q_unbuf <= my_rom(4230);
      when "1000010000111" => q_unbuf <= my_rom(4231);
      when "1000010001000" => q_unbuf <= my_rom(4232);
      when "1000010001001" => q_unbuf <= my_rom(4233);
      when "1000010001010" => q_unbuf <= my_rom(4234);
      when "1000010001011" => q_unbuf <= my_rom(4235);
      when "1000010001100" => q_unbuf <= my_rom(4236);
      when "1000010001101" => q_unbuf <= my_rom(4237);
      when "1000010001110" => q_unbuf <= my_rom(4238);
      when "1000010001111" => q_unbuf <= my_rom(4239);
      when "1000010010000" => q_unbuf <= my_rom(4240);
      when "1000010010001" => q_unbuf <= my_rom(4241);
      when "1000010010010" => q_unbuf <= my_rom(4242);
      when "1000010010011" => q_unbuf <= my_rom(4243);
      when "1000010010100" => q_unbuf <= my_rom(4244);
      when "1000010010101" => q_unbuf <= my_rom(4245);
      when "1000010010110" => q_unbuf <= my_rom(4246);
      when "1000010010111" => q_unbuf <= my_rom(4247);
      when "1000010011000" => q_unbuf <= my_rom(4248);
      when "1000010011001" => q_unbuf <= my_rom(4249);
      when "1000010011010" => q_unbuf <= my_rom(4250);
      when "1000010011011" => q_unbuf <= my_rom(4251);
      when "1000010011100" => q_unbuf <= my_rom(4252);
      when "1000010011101" => q_unbuf <= my_rom(4253);
      when "1000010011110" => q_unbuf <= my_rom(4254);
      when "1000010011111" => q_unbuf <= my_rom(4255);
      when "1000010100000" => q_unbuf <= my_rom(4256);
      when "1000010100001" => q_unbuf <= my_rom(4257);
      when "1000010100010" => q_unbuf <= my_rom(4258);
      when "1000010100011" => q_unbuf <= my_rom(4259);
      when "1000010100100" => q_unbuf <= my_rom(4260);
      when "1000010100101" => q_unbuf <= my_rom(4261);
      when "1000010100110" => q_unbuf <= my_rom(4262);
      when "1000010100111" => q_unbuf <= my_rom(4263);
      when "1000010101000" => q_unbuf <= my_rom(4264);
      when "1000010101001" => q_unbuf <= my_rom(4265);
      when "1000010101010" => q_unbuf <= my_rom(4266);
      when "1000010101011" => q_unbuf <= my_rom(4267);
      when "1000010101100" => q_unbuf <= my_rom(4268);
      when "1000010101101" => q_unbuf <= my_rom(4269);
      when "1000010101110" => q_unbuf <= my_rom(4270);
      when "1000010101111" => q_unbuf <= my_rom(4271);
      when "1000010110000" => q_unbuf <= my_rom(4272);
      when "1000010110001" => q_unbuf <= my_rom(4273);
      when "1000010110010" => q_unbuf <= my_rom(4274);
      when "1000010110011" => q_unbuf <= my_rom(4275);
      when "1000010110100" => q_unbuf <= my_rom(4276);
      when "1000010110101" => q_unbuf <= my_rom(4277);
      when "1000010110110" => q_unbuf <= my_rom(4278);
      when "1000010110111" => q_unbuf <= my_rom(4279);
      when "1000010111000" => q_unbuf <= my_rom(4280);
      when "1000010111001" => q_unbuf <= my_rom(4281);
      when "1000010111010" => q_unbuf <= my_rom(4282);
      when "1000010111011" => q_unbuf <= my_rom(4283);
      when "1000010111100" => q_unbuf <= my_rom(4284);
      when "1000010111101" => q_unbuf <= my_rom(4285);
      when "1000010111110" => q_unbuf <= my_rom(4286);
      when "1000010111111" => q_unbuf <= my_rom(4287);
      when "1000011000000" => q_unbuf <= my_rom(4288);
      when "1000011000001" => q_unbuf <= my_rom(4289);
      when "1000011000010" => q_unbuf <= my_rom(4290);
      when "1000011000011" => q_unbuf <= my_rom(4291);
      when "1000011000100" => q_unbuf <= my_rom(4292);
      when "1000011000101" => q_unbuf <= my_rom(4293);
      when "1000011000110" => q_unbuf <= my_rom(4294);
      when "1000011000111" => q_unbuf <= my_rom(4295);
      when "1000011001000" => q_unbuf <= my_rom(4296);
      when "1000011001001" => q_unbuf <= my_rom(4297);
      when "1000011001010" => q_unbuf <= my_rom(4298);
      when "1000011001011" => q_unbuf <= my_rom(4299);
      when "1000011001100" => q_unbuf <= my_rom(4300);
      when "1000011001101" => q_unbuf <= my_rom(4301);
      when "1000011001110" => q_unbuf <= my_rom(4302);
      when "1000011001111" => q_unbuf <= my_rom(4303);
      when "1000011010000" => q_unbuf <= my_rom(4304);
      when "1000011010001" => q_unbuf <= my_rom(4305);
      when "1000011010010" => q_unbuf <= my_rom(4306);
      when "1000011010011" => q_unbuf <= my_rom(4307);
      when "1000011010100" => q_unbuf <= my_rom(4308);
      when "1000011010101" => q_unbuf <= my_rom(4309);
      when "1000011010110" => q_unbuf <= my_rom(4310);
      when "1000011010111" => q_unbuf <= my_rom(4311);
      when "1000011011000" => q_unbuf <= my_rom(4312);
      when "1000011011001" => q_unbuf <= my_rom(4313);
      when "1000011011010" => q_unbuf <= my_rom(4314);
      when "1000011011011" => q_unbuf <= my_rom(4315);
      when "1000011011100" => q_unbuf <= my_rom(4316);
      when "1000011011101" => q_unbuf <= my_rom(4317);
      when "1000011011110" => q_unbuf <= my_rom(4318);
      when "1000011011111" => q_unbuf <= my_rom(4319);
      when "1000011100000" => q_unbuf <= my_rom(4320);
      when "1000011100001" => q_unbuf <= my_rom(4321);
      when "1000011100010" => q_unbuf <= my_rom(4322);
      when "1000011100011" => q_unbuf <= my_rom(4323);
      when "1000011100100" => q_unbuf <= my_rom(4324);
      when "1000011100101" => q_unbuf <= my_rom(4325);
      when "1000011100110" => q_unbuf <= my_rom(4326);
      when "1000011100111" => q_unbuf <= my_rom(4327);
      when "1000011101000" => q_unbuf <= my_rom(4328);
      when "1000011101001" => q_unbuf <= my_rom(4329);
      when "1000011101010" => q_unbuf <= my_rom(4330);
      when "1000011101011" => q_unbuf <= my_rom(4331);
      when "1000011101100" => q_unbuf <= my_rom(4332);
      when "1000011101101" => q_unbuf <= my_rom(4333);
      when "1000011101110" => q_unbuf <= my_rom(4334);
      when "1000011101111" => q_unbuf <= my_rom(4335);
      when "1000011110000" => q_unbuf <= my_rom(4336);
      when "1000011110001" => q_unbuf <= my_rom(4337);
      when "1000011110010" => q_unbuf <= my_rom(4338);
      when "1000011110011" => q_unbuf <= my_rom(4339);
      when "1000011110100" => q_unbuf <= my_rom(4340);
      when "1000011110101" => q_unbuf <= my_rom(4341);
      when "1000011110110" => q_unbuf <= my_rom(4342);
      when "1000011110111" => q_unbuf <= my_rom(4343);
      when "1000011111000" => q_unbuf <= my_rom(4344);
      when "1000011111001" => q_unbuf <= my_rom(4345);
      when "1000011111010" => q_unbuf <= my_rom(4346);
      when "1000011111011" => q_unbuf <= my_rom(4347);
      when "1000011111100" => q_unbuf <= my_rom(4348);
      when "1000011111101" => q_unbuf <= my_rom(4349);
      when "1000011111110" => q_unbuf <= my_rom(4350);
      when "1000011111111" => q_unbuf <= my_rom(4351);
      when "1000100000000" => q_unbuf <= my_rom(4352);
      when "1000100000001" => q_unbuf <= my_rom(4353);
      when "1000100000010" => q_unbuf <= my_rom(4354);
      when "1000100000011" => q_unbuf <= my_rom(4355);
      when "1000100000100" => q_unbuf <= my_rom(4356);
      when "1000100000101" => q_unbuf <= my_rom(4357);
      when "1000100000110" => q_unbuf <= my_rom(4358);
      when "1000100000111" => q_unbuf <= my_rom(4359);
      when "1000100001000" => q_unbuf <= my_rom(4360);
      when "1000100001001" => q_unbuf <= my_rom(4361);
      when "1000100001010" => q_unbuf <= my_rom(4362);
      when "1000100001011" => q_unbuf <= my_rom(4363);
      when "1000100001100" => q_unbuf <= my_rom(4364);
      when "1000100001101" => q_unbuf <= my_rom(4365);
      when "1000100001110" => q_unbuf <= my_rom(4366);
      when "1000100001111" => q_unbuf <= my_rom(4367);
      when "1000100010000" => q_unbuf <= my_rom(4368);
      when "1000100010001" => q_unbuf <= my_rom(4369);
      when "1000100010010" => q_unbuf <= my_rom(4370);
      when "1000100010011" => q_unbuf <= my_rom(4371);
      when "1000100010100" => q_unbuf <= my_rom(4372);
      when "1000100010101" => q_unbuf <= my_rom(4373);
      when "1000100010110" => q_unbuf <= my_rom(4374);
      when "1000100010111" => q_unbuf <= my_rom(4375);
      when "1000100011000" => q_unbuf <= my_rom(4376);
      when "1000100011001" => q_unbuf <= my_rom(4377);
      when "1000100011010" => q_unbuf <= my_rom(4378);
      when "1000100011011" => q_unbuf <= my_rom(4379);
      when "1000100011100" => q_unbuf <= my_rom(4380);
      when "1000100011101" => q_unbuf <= my_rom(4381);
      when "1000100011110" => q_unbuf <= my_rom(4382);
      when "1000100011111" => q_unbuf <= my_rom(4383);
      when "1000100100000" => q_unbuf <= my_rom(4384);
      when "1000100100001" => q_unbuf <= my_rom(4385);
      when "1000100100010" => q_unbuf <= my_rom(4386);
      when "1000100100011" => q_unbuf <= my_rom(4387);
      when "1000100100100" => q_unbuf <= my_rom(4388);
      when "1000100100101" => q_unbuf <= my_rom(4389);
      when "1000100100110" => q_unbuf <= my_rom(4390);
      when "1000100100111" => q_unbuf <= my_rom(4391);
      when "1000100101000" => q_unbuf <= my_rom(4392);
      when "1000100101001" => q_unbuf <= my_rom(4393);
      when "1000100101010" => q_unbuf <= my_rom(4394);
      when "1000100101011" => q_unbuf <= my_rom(4395);
      when "1000100101100" => q_unbuf <= my_rom(4396);
      when "1000100101101" => q_unbuf <= my_rom(4397);
      when "1000100101110" => q_unbuf <= my_rom(4398);
      when "1000100101111" => q_unbuf <= my_rom(4399);
      when "1000100110000" => q_unbuf <= my_rom(4400);
      when "1000100110001" => q_unbuf <= my_rom(4401);
      when "1000100110010" => q_unbuf <= my_rom(4402);
      when "1000100110011" => q_unbuf <= my_rom(4403);
      when "1000100110100" => q_unbuf <= my_rom(4404);
      when "1000100110101" => q_unbuf <= my_rom(4405);
      when "1000100110110" => q_unbuf <= my_rom(4406);
      when "1000100110111" => q_unbuf <= my_rom(4407);
      when "1000100111000" => q_unbuf <= my_rom(4408);
      when "1000100111001" => q_unbuf <= my_rom(4409);
      when "1000100111010" => q_unbuf <= my_rom(4410);
      when "1000100111011" => q_unbuf <= my_rom(4411);
      when "1000100111100" => q_unbuf <= my_rom(4412);
      when "1000100111101" => q_unbuf <= my_rom(4413);
      when "1000100111110" => q_unbuf <= my_rom(4414);
      when "1000100111111" => q_unbuf <= my_rom(4415);
      when "1000101000000" => q_unbuf <= my_rom(4416);
      when "1000101000001" => q_unbuf <= my_rom(4417);
      when "1000101000010" => q_unbuf <= my_rom(4418);
      when "1000101000011" => q_unbuf <= my_rom(4419);
      when "1000101000100" => q_unbuf <= my_rom(4420);
      when "1000101000101" => q_unbuf <= my_rom(4421);
      when "1000101000110" => q_unbuf <= my_rom(4422);
      when "1000101000111" => q_unbuf <= my_rom(4423);
      when "1000101001000" => q_unbuf <= my_rom(4424);
      when "1000101001001" => q_unbuf <= my_rom(4425);
      when "1000101001010" => q_unbuf <= my_rom(4426);
      when "1000101001011" => q_unbuf <= my_rom(4427);
      when "1000101001100" => q_unbuf <= my_rom(4428);
      when "1000101001101" => q_unbuf <= my_rom(4429);
      when "1000101001110" => q_unbuf <= my_rom(4430);
      when "1000101001111" => q_unbuf <= my_rom(4431);
      when "1000101010000" => q_unbuf <= my_rom(4432);
      when "1000101010001" => q_unbuf <= my_rom(4433);
      when "1000101010010" => q_unbuf <= my_rom(4434);
      when "1000101010011" => q_unbuf <= my_rom(4435);
      when "1000101010100" => q_unbuf <= my_rom(4436);
      when "1000101010101" => q_unbuf <= my_rom(4437);
      when "1000101010110" => q_unbuf <= my_rom(4438);
      when "1000101010111" => q_unbuf <= my_rom(4439);
      when "1000101011000" => q_unbuf <= my_rom(4440);
      when "1000101011001" => q_unbuf <= my_rom(4441);
      when "1000101011010" => q_unbuf <= my_rom(4442);
      when "1000101011011" => q_unbuf <= my_rom(4443);
      when "1000101011100" => q_unbuf <= my_rom(4444);
      when "1000101011101" => q_unbuf <= my_rom(4445);
      when "1000101011110" => q_unbuf <= my_rom(4446);
      when "1000101011111" => q_unbuf <= my_rom(4447);
      when "1000101100000" => q_unbuf <= my_rom(4448);
      when "1000101100001" => q_unbuf <= my_rom(4449);
      when "1000101100010" => q_unbuf <= my_rom(4450);
      when "1000101100011" => q_unbuf <= my_rom(4451);
      when "1000101100100" => q_unbuf <= my_rom(4452);
      when "1000101100101" => q_unbuf <= my_rom(4453);
      when "1000101100110" => q_unbuf <= my_rom(4454);
      when "1000101100111" => q_unbuf <= my_rom(4455);
      when "1000101101000" => q_unbuf <= my_rom(4456);
      when "1000101101001" => q_unbuf <= my_rom(4457);
      when "1000101101010" => q_unbuf <= my_rom(4458);
      when "1000101101011" => q_unbuf <= my_rom(4459);
      when "1000101101100" => q_unbuf <= my_rom(4460);
      when "1000101101101" => q_unbuf <= my_rom(4461);
      when "1000101101110" => q_unbuf <= my_rom(4462);
      when "1000101101111" => q_unbuf <= my_rom(4463);
      when "1000101110000" => q_unbuf <= my_rom(4464);
      when "1000101110001" => q_unbuf <= my_rom(4465);
      when "1000101110010" => q_unbuf <= my_rom(4466);
      when "1000101110011" => q_unbuf <= my_rom(4467);
      when "1000101110100" => q_unbuf <= my_rom(4468);
      when "1000101110101" => q_unbuf <= my_rom(4469);
      when "1000101110110" => q_unbuf <= my_rom(4470);
      when "1000101110111" => q_unbuf <= my_rom(4471);
      when "1000101111000" => q_unbuf <= my_rom(4472);
      when "1000101111001" => q_unbuf <= my_rom(4473);
      when "1000101111010" => q_unbuf <= my_rom(4474);
      when "1000101111011" => q_unbuf <= my_rom(4475);
      when "1000101111100" => q_unbuf <= my_rom(4476);
      when "1000101111101" => q_unbuf <= my_rom(4477);
      when "1000101111110" => q_unbuf <= my_rom(4478);
      when "1000101111111" => q_unbuf <= my_rom(4479);
      when "1000110000000" => q_unbuf <= my_rom(4480);
      when "1000110000001" => q_unbuf <= my_rom(4481);
      when "1000110000010" => q_unbuf <= my_rom(4482);
      when "1000110000011" => q_unbuf <= my_rom(4483);
      when "1000110000100" => q_unbuf <= my_rom(4484);
      when "1000110000101" => q_unbuf <= my_rom(4485);
      when "1000110000110" => q_unbuf <= my_rom(4486);
      when "1000110000111" => q_unbuf <= my_rom(4487);
      when "1000110001000" => q_unbuf <= my_rom(4488);
      when "1000110001001" => q_unbuf <= my_rom(4489);
      when "1000110001010" => q_unbuf <= my_rom(4490);
      when "1000110001011" => q_unbuf <= my_rom(4491);
      when "1000110001100" => q_unbuf <= my_rom(4492);
      when "1000110001101" => q_unbuf <= my_rom(4493);
      when "1000110001110" => q_unbuf <= my_rom(4494);
      when "1000110001111" => q_unbuf <= my_rom(4495);
      when "1000110010000" => q_unbuf <= my_rom(4496);
      when "1000110010001" => q_unbuf <= my_rom(4497);
      when "1000110010010" => q_unbuf <= my_rom(4498);
      when "1000110010011" => q_unbuf <= my_rom(4499);
      when "1000110010100" => q_unbuf <= my_rom(4500);
      when "1000110010101" => q_unbuf <= my_rom(4501);
      when "1000110010110" => q_unbuf <= my_rom(4502);
      when "1000110010111" => q_unbuf <= my_rom(4503);
      when "1000110011000" => q_unbuf <= my_rom(4504);
      when "1000110011001" => q_unbuf <= my_rom(4505);
      when "1000110011010" => q_unbuf <= my_rom(4506);
      when "1000110011011" => q_unbuf <= my_rom(4507);
      when "1000110011100" => q_unbuf <= my_rom(4508);
      when "1000110011101" => q_unbuf <= my_rom(4509);
      when "1000110011110" => q_unbuf <= my_rom(4510);
      when "1000110011111" => q_unbuf <= my_rom(4511);
      when "1000110100000" => q_unbuf <= my_rom(4512);
      when "1000110100001" => q_unbuf <= my_rom(4513);
      when "1000110100010" => q_unbuf <= my_rom(4514);
      when "1000110100011" => q_unbuf <= my_rom(4515);
      when "1000110100100" => q_unbuf <= my_rom(4516);
      when "1000110100101" => q_unbuf <= my_rom(4517);
      when "1000110100110" => q_unbuf <= my_rom(4518);
      when "1000110100111" => q_unbuf <= my_rom(4519);
      when "1000110101000" => q_unbuf <= my_rom(4520);
      when "1000110101001" => q_unbuf <= my_rom(4521);
      when "1000110101010" => q_unbuf <= my_rom(4522);
      when "1000110101011" => q_unbuf <= my_rom(4523);
      when "1000110101100" => q_unbuf <= my_rom(4524);
      when "1000110101101" => q_unbuf <= my_rom(4525);
      when "1000110101110" => q_unbuf <= my_rom(4526);
      when "1000110101111" => q_unbuf <= my_rom(4527);
      when "1000110110000" => q_unbuf <= my_rom(4528);
      when "1000110110001" => q_unbuf <= my_rom(4529);
      when "1000110110010" => q_unbuf <= my_rom(4530);
      when "1000110110011" => q_unbuf <= my_rom(4531);
      when "1000110110100" => q_unbuf <= my_rom(4532);
      when "1000110110101" => q_unbuf <= my_rom(4533);
      when "1000110110110" => q_unbuf <= my_rom(4534);
      when "1000110110111" => q_unbuf <= my_rom(4535);
      when "1000110111000" => q_unbuf <= my_rom(4536);
      when "1000110111001" => q_unbuf <= my_rom(4537);
      when "1000110111010" => q_unbuf <= my_rom(4538);
      when "1000110111011" => q_unbuf <= my_rom(4539);
      when "1000110111100" => q_unbuf <= my_rom(4540);
      when "1000110111101" => q_unbuf <= my_rom(4541);
      when "1000110111110" => q_unbuf <= my_rom(4542);
      when "1000110111111" => q_unbuf <= my_rom(4543);
      when "1000111000000" => q_unbuf <= my_rom(4544);
      when "1000111000001" => q_unbuf <= my_rom(4545);
      when "1000111000010" => q_unbuf <= my_rom(4546);
      when "1000111000011" => q_unbuf <= my_rom(4547);
      when "1000111000100" => q_unbuf <= my_rom(4548);
      when "1000111000101" => q_unbuf <= my_rom(4549);
      when "1000111000110" => q_unbuf <= my_rom(4550);
      when "1000111000111" => q_unbuf <= my_rom(4551);
      when "1000111001000" => q_unbuf <= my_rom(4552);
      when "1000111001001" => q_unbuf <= my_rom(4553);
      when "1000111001010" => q_unbuf <= my_rom(4554);
      when "1000111001011" => q_unbuf <= my_rom(4555);
      when "1000111001100" => q_unbuf <= my_rom(4556);
      when "1000111001101" => q_unbuf <= my_rom(4557);
      when "1000111001110" => q_unbuf <= my_rom(4558);
      when "1000111001111" => q_unbuf <= my_rom(4559);
      when "1000111010000" => q_unbuf <= my_rom(4560);
      when "1000111010001" => q_unbuf <= my_rom(4561);
      when "1000111010010" => q_unbuf <= my_rom(4562);
      when "1000111010011" => q_unbuf <= my_rom(4563);
      when "1000111010100" => q_unbuf <= my_rom(4564);
      when "1000111010101" => q_unbuf <= my_rom(4565);
      when "1000111010110" => q_unbuf <= my_rom(4566);
      when "1000111010111" => q_unbuf <= my_rom(4567);
      when "1000111011000" => q_unbuf <= my_rom(4568);
      when "1000111011001" => q_unbuf <= my_rom(4569);
      when "1000111011010" => q_unbuf <= my_rom(4570);
      when "1000111011011" => q_unbuf <= my_rom(4571);
      when "1000111011100" => q_unbuf <= my_rom(4572);
      when "1000111011101" => q_unbuf <= my_rom(4573);
      when "1000111011110" => q_unbuf <= my_rom(4574);
      when "1000111011111" => q_unbuf <= my_rom(4575);
      when "1000111100000" => q_unbuf <= my_rom(4576);
      when "1000111100001" => q_unbuf <= my_rom(4577);
      when "1000111100010" => q_unbuf <= my_rom(4578);
      when "1000111100011" => q_unbuf <= my_rom(4579);
      when "1000111100100" => q_unbuf <= my_rom(4580);
      when "1000111100101" => q_unbuf <= my_rom(4581);
      when "1000111100110" => q_unbuf <= my_rom(4582);
      when "1000111100111" => q_unbuf <= my_rom(4583);
      when "1000111101000" => q_unbuf <= my_rom(4584);
      when "1000111101001" => q_unbuf <= my_rom(4585);
      when "1000111101010" => q_unbuf <= my_rom(4586);
      when "1000111101011" => q_unbuf <= my_rom(4587);
      when "1000111101100" => q_unbuf <= my_rom(4588);
      when "1000111101101" => q_unbuf <= my_rom(4589);
      when "1000111101110" => q_unbuf <= my_rom(4590);
      when "1000111101111" => q_unbuf <= my_rom(4591);
      when "1000111110000" => q_unbuf <= my_rom(4592);
      when "1000111110001" => q_unbuf <= my_rom(4593);
      when "1000111110010" => q_unbuf <= my_rom(4594);
      when "1000111110011" => q_unbuf <= my_rom(4595);
      when "1000111110100" => q_unbuf <= my_rom(4596);
      when "1000111110101" => q_unbuf <= my_rom(4597);
      when "1000111110110" => q_unbuf <= my_rom(4598);
      when "1000111110111" => q_unbuf <= my_rom(4599);
      when "1000111111000" => q_unbuf <= my_rom(4600);
      when "1000111111001" => q_unbuf <= my_rom(4601);
      when "1000111111010" => q_unbuf <= my_rom(4602);
      when "1000111111011" => q_unbuf <= my_rom(4603);
      when "1000111111100" => q_unbuf <= my_rom(4604);
      when "1000111111101" => q_unbuf <= my_rom(4605);
      when "1000111111110" => q_unbuf <= my_rom(4606);
      when "1000111111111" => q_unbuf <= my_rom(4607);
      when "1001000000000" => q_unbuf <= my_rom(4608);
      when "1001000000001" => q_unbuf <= my_rom(4609);
      when "1001000000010" => q_unbuf <= my_rom(4610);
      when "1001000000011" => q_unbuf <= my_rom(4611);
      when "1001000000100" => q_unbuf <= my_rom(4612);
      when "1001000000101" => q_unbuf <= my_rom(4613);
      when "1001000000110" => q_unbuf <= my_rom(4614);
      when "1001000000111" => q_unbuf <= my_rom(4615);
      when "1001000001000" => q_unbuf <= my_rom(4616);
      when "1001000001001" => q_unbuf <= my_rom(4617);
      when "1001000001010" => q_unbuf <= my_rom(4618);
      when "1001000001011" => q_unbuf <= my_rom(4619);
      when "1001000001100" => q_unbuf <= my_rom(4620);
      when "1001000001101" => q_unbuf <= my_rom(4621);
      when "1001000001110" => q_unbuf <= my_rom(4622);
      when "1001000001111" => q_unbuf <= my_rom(4623);
      when "1001000010000" => q_unbuf <= my_rom(4624);
      when "1001000010001" => q_unbuf <= my_rom(4625);
      when "1001000010010" => q_unbuf <= my_rom(4626);
      when "1001000010011" => q_unbuf <= my_rom(4627);
      when "1001000010100" => q_unbuf <= my_rom(4628);
      when "1001000010101" => q_unbuf <= my_rom(4629);
      when "1001000010110" => q_unbuf <= my_rom(4630);
      when "1001000010111" => q_unbuf <= my_rom(4631);
      when "1001000011000" => q_unbuf <= my_rom(4632);
      when "1001000011001" => q_unbuf <= my_rom(4633);
      when "1001000011010" => q_unbuf <= my_rom(4634);
      when "1001000011011" => q_unbuf <= my_rom(4635);
      when "1001000011100" => q_unbuf <= my_rom(4636);
      when "1001000011101" => q_unbuf <= my_rom(4637);
      when "1001000011110" => q_unbuf <= my_rom(4638);
      when "1001000011111" => q_unbuf <= my_rom(4639);
      when "1001000100000" => q_unbuf <= my_rom(4640);
      when "1001000100001" => q_unbuf <= my_rom(4641);
      when "1001000100010" => q_unbuf <= my_rom(4642);
      when "1001000100011" => q_unbuf <= my_rom(4643);
      when "1001000100100" => q_unbuf <= my_rom(4644);
      when "1001000100101" => q_unbuf <= my_rom(4645);
      when "1001000100110" => q_unbuf <= my_rom(4646);
      when "1001000100111" => q_unbuf <= my_rom(4647);
      when "1001000101000" => q_unbuf <= my_rom(4648);
      when "1001000101001" => q_unbuf <= my_rom(4649);
      when "1001000101010" => q_unbuf <= my_rom(4650);
      when "1001000101011" => q_unbuf <= my_rom(4651);
      when "1001000101100" => q_unbuf <= my_rom(4652);
      when "1001000101101" => q_unbuf <= my_rom(4653);
      when "1001000101110" => q_unbuf <= my_rom(4654);
      when "1001000101111" => q_unbuf <= my_rom(4655);
      when "1001000110000" => q_unbuf <= my_rom(4656);
      when "1001000110001" => q_unbuf <= my_rom(4657);
      when "1001000110010" => q_unbuf <= my_rom(4658);
      when "1001000110011" => q_unbuf <= my_rom(4659);
      when "1001000110100" => q_unbuf <= my_rom(4660);
      when "1001000110101" => q_unbuf <= my_rom(4661);
      when "1001000110110" => q_unbuf <= my_rom(4662);
      when "1001000110111" => q_unbuf <= my_rom(4663);
      when "1001000111000" => q_unbuf <= my_rom(4664);
      when "1001000111001" => q_unbuf <= my_rom(4665);
      when "1001000111010" => q_unbuf <= my_rom(4666);
      when "1001000111011" => q_unbuf <= my_rom(4667);
      when "1001000111100" => q_unbuf <= my_rom(4668);
      when "1001000111101" => q_unbuf <= my_rom(4669);
      when "1001000111110" => q_unbuf <= my_rom(4670);
      when "1001000111111" => q_unbuf <= my_rom(4671);
      when "1001001000000" => q_unbuf <= my_rom(4672);
      when "1001001000001" => q_unbuf <= my_rom(4673);
      when "1001001000010" => q_unbuf <= my_rom(4674);
      when "1001001000011" => q_unbuf <= my_rom(4675);
      when "1001001000100" => q_unbuf <= my_rom(4676);
      when "1001001000101" => q_unbuf <= my_rom(4677);
      when "1001001000110" => q_unbuf <= my_rom(4678);
      when "1001001000111" => q_unbuf <= my_rom(4679);
      when "1001001001000" => q_unbuf <= my_rom(4680);
      when "1001001001001" => q_unbuf <= my_rom(4681);
      when "1001001001010" => q_unbuf <= my_rom(4682);
      when "1001001001011" => q_unbuf <= my_rom(4683);
      when "1001001001100" => q_unbuf <= my_rom(4684);
      when "1001001001101" => q_unbuf <= my_rom(4685);
      when "1001001001110" => q_unbuf <= my_rom(4686);
      when "1001001001111" => q_unbuf <= my_rom(4687);
      when "1001001010000" => q_unbuf <= my_rom(4688);
      when "1001001010001" => q_unbuf <= my_rom(4689);
      when "1001001010010" => q_unbuf <= my_rom(4690);
      when "1001001010011" => q_unbuf <= my_rom(4691);
      when "1001001010100" => q_unbuf <= my_rom(4692);
      when "1001001010101" => q_unbuf <= my_rom(4693);
      when "1001001010110" => q_unbuf <= my_rom(4694);
      when "1001001010111" => q_unbuf <= my_rom(4695);
      when "1001001011000" => q_unbuf <= my_rom(4696);
      when "1001001011001" => q_unbuf <= my_rom(4697);
      when "1001001011010" => q_unbuf <= my_rom(4698);
      when "1001001011011" => q_unbuf <= my_rom(4699);
      when "1001001011100" => q_unbuf <= my_rom(4700);
      when "1001001011101" => q_unbuf <= my_rom(4701);
      when "1001001011110" => q_unbuf <= my_rom(4702);
      when "1001001011111" => q_unbuf <= my_rom(4703);
      when "1001001100000" => q_unbuf <= my_rom(4704);
      when "1001001100001" => q_unbuf <= my_rom(4705);
      when "1001001100010" => q_unbuf <= my_rom(4706);
      when "1001001100011" => q_unbuf <= my_rom(4707);
      when "1001001100100" => q_unbuf <= my_rom(4708);
      when "1001001100101" => q_unbuf <= my_rom(4709);
      when "1001001100110" => q_unbuf <= my_rom(4710);
      when "1001001100111" => q_unbuf <= my_rom(4711);
      when "1001001101000" => q_unbuf <= my_rom(4712);
      when "1001001101001" => q_unbuf <= my_rom(4713);
      when "1001001101010" => q_unbuf <= my_rom(4714);
      when "1001001101011" => q_unbuf <= my_rom(4715);
      when "1001001101100" => q_unbuf <= my_rom(4716);
      when "1001001101101" => q_unbuf <= my_rom(4717);
      when "1001001101110" => q_unbuf <= my_rom(4718);
      when "1001001101111" => q_unbuf <= my_rom(4719);
      when "1001001110000" => q_unbuf <= my_rom(4720);
      when "1001001110001" => q_unbuf <= my_rom(4721);
      when "1001001110010" => q_unbuf <= my_rom(4722);
      when "1001001110011" => q_unbuf <= my_rom(4723);
      when "1001001110100" => q_unbuf <= my_rom(4724);
      when "1001001110101" => q_unbuf <= my_rom(4725);
      when "1001001110110" => q_unbuf <= my_rom(4726);
      when "1001001110111" => q_unbuf <= my_rom(4727);
      when "1001001111000" => q_unbuf <= my_rom(4728);
      when "1001001111001" => q_unbuf <= my_rom(4729);
      when "1001001111010" => q_unbuf <= my_rom(4730);
      when "1001001111011" => q_unbuf <= my_rom(4731);
      when "1001001111100" => q_unbuf <= my_rom(4732);
      when "1001001111101" => q_unbuf <= my_rom(4733);
      when "1001001111110" => q_unbuf <= my_rom(4734);
      when "1001001111111" => q_unbuf <= my_rom(4735);
      when "1001010000000" => q_unbuf <= my_rom(4736);
      when "1001010000001" => q_unbuf <= my_rom(4737);
      when "1001010000010" => q_unbuf <= my_rom(4738);
      when "1001010000011" => q_unbuf <= my_rom(4739);
      when "1001010000100" => q_unbuf <= my_rom(4740);
      when "1001010000101" => q_unbuf <= my_rom(4741);
      when "1001010000110" => q_unbuf <= my_rom(4742);
      when "1001010000111" => q_unbuf <= my_rom(4743);
      when "1001010001000" => q_unbuf <= my_rom(4744);
      when "1001010001001" => q_unbuf <= my_rom(4745);
      when "1001010001010" => q_unbuf <= my_rom(4746);
      when "1001010001011" => q_unbuf <= my_rom(4747);
      when "1001010001100" => q_unbuf <= my_rom(4748);
      when "1001010001101" => q_unbuf <= my_rom(4749);
      when "1001010001110" => q_unbuf <= my_rom(4750);
      when "1001010001111" => q_unbuf <= my_rom(4751);
      when "1001010010000" => q_unbuf <= my_rom(4752);
      when "1001010010001" => q_unbuf <= my_rom(4753);
      when "1001010010010" => q_unbuf <= my_rom(4754);
      when "1001010010011" => q_unbuf <= my_rom(4755);
      when "1001010010100" => q_unbuf <= my_rom(4756);
      when "1001010010101" => q_unbuf <= my_rom(4757);
      when "1001010010110" => q_unbuf <= my_rom(4758);
      when "1001010010111" => q_unbuf <= my_rom(4759);
      when "1001010011000" => q_unbuf <= my_rom(4760);
      when "1001010011001" => q_unbuf <= my_rom(4761);
      when "1001010011010" => q_unbuf <= my_rom(4762);
      when "1001010011011" => q_unbuf <= my_rom(4763);
      when "1001010011100" => q_unbuf <= my_rom(4764);
      when "1001010011101" => q_unbuf <= my_rom(4765);
      when "1001010011110" => q_unbuf <= my_rom(4766);
      when "1001010011111" => q_unbuf <= my_rom(4767);
      when "1001010100000" => q_unbuf <= my_rom(4768);
      when "1001010100001" => q_unbuf <= my_rom(4769);
      when "1001010100010" => q_unbuf <= my_rom(4770);
      when "1001010100011" => q_unbuf <= my_rom(4771);
      when "1001010100100" => q_unbuf <= my_rom(4772);
      when "1001010100101" => q_unbuf <= my_rom(4773);
      when "1001010100110" => q_unbuf <= my_rom(4774);
      when "1001010100111" => q_unbuf <= my_rom(4775);
      when "1001010101000" => q_unbuf <= my_rom(4776);
      when "1001010101001" => q_unbuf <= my_rom(4777);
      when "1001010101010" => q_unbuf <= my_rom(4778);
      when "1001010101011" => q_unbuf <= my_rom(4779);
      when "1001010101100" => q_unbuf <= my_rom(4780);
      when "1001010101101" => q_unbuf <= my_rom(4781);
      when "1001010101110" => q_unbuf <= my_rom(4782);
      when "1001010101111" => q_unbuf <= my_rom(4783);
      when "1001010110000" => q_unbuf <= my_rom(4784);
      when "1001010110001" => q_unbuf <= my_rom(4785);
      when "1001010110010" => q_unbuf <= my_rom(4786);
      when "1001010110011" => q_unbuf <= my_rom(4787);
      when "1001010110100" => q_unbuf <= my_rom(4788);
      when "1001010110101" => q_unbuf <= my_rom(4789);
      when "1001010110110" => q_unbuf <= my_rom(4790);
      when "1001010110111" => q_unbuf <= my_rom(4791);
      when "1001010111000" => q_unbuf <= my_rom(4792);
      when "1001010111001" => q_unbuf <= my_rom(4793);
      when "1001010111010" => q_unbuf <= my_rom(4794);
      when "1001010111011" => q_unbuf <= my_rom(4795);
      when "1001010111100" => q_unbuf <= my_rom(4796);
      when "1001010111101" => q_unbuf <= my_rom(4797);
      when "1001010111110" => q_unbuf <= my_rom(4798);
      when "1001010111111" => q_unbuf <= my_rom(4799);
      when "1001011000000" => q_unbuf <= my_rom(4800);
      when "1001011000001" => q_unbuf <= my_rom(4801);
      when "1001011000010" => q_unbuf <= my_rom(4802);
      when "1001011000011" => q_unbuf <= my_rom(4803);
      when "1001011000100" => q_unbuf <= my_rom(4804);
      when "1001011000101" => q_unbuf <= my_rom(4805);
      when "1001011000110" => q_unbuf <= my_rom(4806);
      when "1001011000111" => q_unbuf <= my_rom(4807);
      when "1001011001000" => q_unbuf <= my_rom(4808);
      when "1001011001001" => q_unbuf <= my_rom(4809);
      when "1001011001010" => q_unbuf <= my_rom(4810);
      when "1001011001011" => q_unbuf <= my_rom(4811);
      when "1001011001100" => q_unbuf <= my_rom(4812);
      when "1001011001101" => q_unbuf <= my_rom(4813);
      when "1001011001110" => q_unbuf <= my_rom(4814);
      when "1001011001111" => q_unbuf <= my_rom(4815);
      when "1001011010000" => q_unbuf <= my_rom(4816);
      when "1001011010001" => q_unbuf <= my_rom(4817);
      when "1001011010010" => q_unbuf <= my_rom(4818);
      when "1001011010011" => q_unbuf <= my_rom(4819);
      when "1001011010100" => q_unbuf <= my_rom(4820);
      when "1001011010101" => q_unbuf <= my_rom(4821);
      when "1001011010110" => q_unbuf <= my_rom(4822);
      when "1001011010111" => q_unbuf <= my_rom(4823);
      when "1001011011000" => q_unbuf <= my_rom(4824);
      when "1001011011001" => q_unbuf <= my_rom(4825);
      when "1001011011010" => q_unbuf <= my_rom(4826);
      when "1001011011011" => q_unbuf <= my_rom(4827);
      when "1001011011100" => q_unbuf <= my_rom(4828);
      when "1001011011101" => q_unbuf <= my_rom(4829);
      when "1001011011110" => q_unbuf <= my_rom(4830);
      when "1001011011111" => q_unbuf <= my_rom(4831);
      when "1001011100000" => q_unbuf <= my_rom(4832);
      when "1001011100001" => q_unbuf <= my_rom(4833);
      when "1001011100010" => q_unbuf <= my_rom(4834);
      when "1001011100011" => q_unbuf <= my_rom(4835);
      when "1001011100100" => q_unbuf <= my_rom(4836);
      when "1001011100101" => q_unbuf <= my_rom(4837);
      when "1001011100110" => q_unbuf <= my_rom(4838);
      when "1001011100111" => q_unbuf <= my_rom(4839);
      when "1001011101000" => q_unbuf <= my_rom(4840);
      when "1001011101001" => q_unbuf <= my_rom(4841);
      when "1001011101010" => q_unbuf <= my_rom(4842);
      when "1001011101011" => q_unbuf <= my_rom(4843);
      when "1001011101100" => q_unbuf <= my_rom(4844);
      when "1001011101101" => q_unbuf <= my_rom(4845);
      when "1001011101110" => q_unbuf <= my_rom(4846);
      when "1001011101111" => q_unbuf <= my_rom(4847);
      when "1001011110000" => q_unbuf <= my_rom(4848);
      when "1001011110001" => q_unbuf <= my_rom(4849);
      when "1001011110010" => q_unbuf <= my_rom(4850);
      when "1001011110011" => q_unbuf <= my_rom(4851);
      when "1001011110100" => q_unbuf <= my_rom(4852);
      when "1001011110101" => q_unbuf <= my_rom(4853);
      when "1001011110110" => q_unbuf <= my_rom(4854);
      when "1001011110111" => q_unbuf <= my_rom(4855);
      when "1001011111000" => q_unbuf <= my_rom(4856);
      when "1001011111001" => q_unbuf <= my_rom(4857);
      when "1001011111010" => q_unbuf <= my_rom(4858);
      when "1001011111011" => q_unbuf <= my_rom(4859);
      when "1001011111100" => q_unbuf <= my_rom(4860);
      when "1001011111101" => q_unbuf <= my_rom(4861);
      when "1001011111110" => q_unbuf <= my_rom(4862);
      when "1001011111111" => q_unbuf <= my_rom(4863);
      when "1001100000000" => q_unbuf <= my_rom(4864);
      when "1001100000001" => q_unbuf <= my_rom(4865);
      when "1001100000010" => q_unbuf <= my_rom(4866);
      when "1001100000011" => q_unbuf <= my_rom(4867);
      when "1001100000100" => q_unbuf <= my_rom(4868);
      when "1001100000101" => q_unbuf <= my_rom(4869);
      when "1001100000110" => q_unbuf <= my_rom(4870);
      when "1001100000111" => q_unbuf <= my_rom(4871);
      when "1001100001000" => q_unbuf <= my_rom(4872);
      when "1001100001001" => q_unbuf <= my_rom(4873);
      when "1001100001010" => q_unbuf <= my_rom(4874);
      when "1001100001011" => q_unbuf <= my_rom(4875);
      when "1001100001100" => q_unbuf <= my_rom(4876);
      when "1001100001101" => q_unbuf <= my_rom(4877);
      when "1001100001110" => q_unbuf <= my_rom(4878);
      when "1001100001111" => q_unbuf <= my_rom(4879);
      when "1001100010000" => q_unbuf <= my_rom(4880);
      when "1001100010001" => q_unbuf <= my_rom(4881);
      when "1001100010010" => q_unbuf <= my_rom(4882);
      when "1001100010011" => q_unbuf <= my_rom(4883);
      when "1001100010100" => q_unbuf <= my_rom(4884);
      when "1001100010101" => q_unbuf <= my_rom(4885);
      when "1001100010110" => q_unbuf <= my_rom(4886);
      when "1001100010111" => q_unbuf <= my_rom(4887);
      when "1001100011000" => q_unbuf <= my_rom(4888);
      when "1001100011001" => q_unbuf <= my_rom(4889);
      when "1001100011010" => q_unbuf <= my_rom(4890);
      when "1001100011011" => q_unbuf <= my_rom(4891);
      when "1001100011100" => q_unbuf <= my_rom(4892);
      when "1001100011101" => q_unbuf <= my_rom(4893);
      when "1001100011110" => q_unbuf <= my_rom(4894);
      when "1001100011111" => q_unbuf <= my_rom(4895);
      when "1001100100000" => q_unbuf <= my_rom(4896);
      when "1001100100001" => q_unbuf <= my_rom(4897);
      when "1001100100010" => q_unbuf <= my_rom(4898);
      when "1001100100011" => q_unbuf <= my_rom(4899);
      when "1001100100100" => q_unbuf <= my_rom(4900);
      when "1001100100101" => q_unbuf <= my_rom(4901);
      when "1001100100110" => q_unbuf <= my_rom(4902);
      when "1001100100111" => q_unbuf <= my_rom(4903);
      when "1001100101000" => q_unbuf <= my_rom(4904);
      when "1001100101001" => q_unbuf <= my_rom(4905);
      when "1001100101010" => q_unbuf <= my_rom(4906);
      when "1001100101011" => q_unbuf <= my_rom(4907);
      when "1001100101100" => q_unbuf <= my_rom(4908);
      when "1001100101101" => q_unbuf <= my_rom(4909);
      when "1001100101110" => q_unbuf <= my_rom(4910);
      when "1001100101111" => q_unbuf <= my_rom(4911);
      when "1001100110000" => q_unbuf <= my_rom(4912);
      when "1001100110001" => q_unbuf <= my_rom(4913);
      when "1001100110010" => q_unbuf <= my_rom(4914);
      when "1001100110011" => q_unbuf <= my_rom(4915);
      when "1001100110100" => q_unbuf <= my_rom(4916);
      when "1001100110101" => q_unbuf <= my_rom(4917);
      when "1001100110110" => q_unbuf <= my_rom(4918);
      when "1001100110111" => q_unbuf <= my_rom(4919);
      when "1001100111000" => q_unbuf <= my_rom(4920);
      when "1001100111001" => q_unbuf <= my_rom(4921);
      when "1001100111010" => q_unbuf <= my_rom(4922);
      when "1001100111011" => q_unbuf <= my_rom(4923);
      when "1001100111100" => q_unbuf <= my_rom(4924);
      when "1001100111101" => q_unbuf <= my_rom(4925);
      when "1001100111110" => q_unbuf <= my_rom(4926);
      when "1001100111111" => q_unbuf <= my_rom(4927);
      when "1001101000000" => q_unbuf <= my_rom(4928);
      when "1001101000001" => q_unbuf <= my_rom(4929);
      when "1001101000010" => q_unbuf <= my_rom(4930);
      when "1001101000011" => q_unbuf <= my_rom(4931);
      when "1001101000100" => q_unbuf <= my_rom(4932);
      when "1001101000101" => q_unbuf <= my_rom(4933);
      when "1001101000110" => q_unbuf <= my_rom(4934);
      when "1001101000111" => q_unbuf <= my_rom(4935);
      when "1001101001000" => q_unbuf <= my_rom(4936);
      when "1001101001001" => q_unbuf <= my_rom(4937);
      when "1001101001010" => q_unbuf <= my_rom(4938);
      when "1001101001011" => q_unbuf <= my_rom(4939);
      when "1001101001100" => q_unbuf <= my_rom(4940);
      when "1001101001101" => q_unbuf <= my_rom(4941);
      when "1001101001110" => q_unbuf <= my_rom(4942);
      when "1001101001111" => q_unbuf <= my_rom(4943);
      when "1001101010000" => q_unbuf <= my_rom(4944);
      when "1001101010001" => q_unbuf <= my_rom(4945);
      when "1001101010010" => q_unbuf <= my_rom(4946);
      when "1001101010011" => q_unbuf <= my_rom(4947);
      when "1001101010100" => q_unbuf <= my_rom(4948);
      when "1001101010101" => q_unbuf <= my_rom(4949);
      when "1001101010110" => q_unbuf <= my_rom(4950);
      when "1001101010111" => q_unbuf <= my_rom(4951);
      when "1001101011000" => q_unbuf <= my_rom(4952);
      when "1001101011001" => q_unbuf <= my_rom(4953);
      when "1001101011010" => q_unbuf <= my_rom(4954);
      when "1001101011011" => q_unbuf <= my_rom(4955);
      when "1001101011100" => q_unbuf <= my_rom(4956);
      when "1001101011101" => q_unbuf <= my_rom(4957);
      when "1001101011110" => q_unbuf <= my_rom(4958);
      when "1001101011111" => q_unbuf <= my_rom(4959);
      when "1001101100000" => q_unbuf <= my_rom(4960);
      when "1001101100001" => q_unbuf <= my_rom(4961);
      when "1001101100010" => q_unbuf <= my_rom(4962);
      when "1001101100011" => q_unbuf <= my_rom(4963);
      when "1001101100100" => q_unbuf <= my_rom(4964);
      when "1001101100101" => q_unbuf <= my_rom(4965);
      when "1001101100110" => q_unbuf <= my_rom(4966);
      when "1001101100111" => q_unbuf <= my_rom(4967);
      when "1001101101000" => q_unbuf <= my_rom(4968);
      when "1001101101001" => q_unbuf <= my_rom(4969);
      when "1001101101010" => q_unbuf <= my_rom(4970);
      when "1001101101011" => q_unbuf <= my_rom(4971);
      when "1001101101100" => q_unbuf <= my_rom(4972);
      when "1001101101101" => q_unbuf <= my_rom(4973);
      when "1001101101110" => q_unbuf <= my_rom(4974);
      when "1001101101111" => q_unbuf <= my_rom(4975);
      when "1001101110000" => q_unbuf <= my_rom(4976);
      when "1001101110001" => q_unbuf <= my_rom(4977);
      when "1001101110010" => q_unbuf <= my_rom(4978);
      when "1001101110011" => q_unbuf <= my_rom(4979);
      when "1001101110100" => q_unbuf <= my_rom(4980);
      when "1001101110101" => q_unbuf <= my_rom(4981);
      when "1001101110110" => q_unbuf <= my_rom(4982);
      when "1001101110111" => q_unbuf <= my_rom(4983);
      when "1001101111000" => q_unbuf <= my_rom(4984);
      when "1001101111001" => q_unbuf <= my_rom(4985);
      when "1001101111010" => q_unbuf <= my_rom(4986);
      when "1001101111011" => q_unbuf <= my_rom(4987);
      when "1001101111100" => q_unbuf <= my_rom(4988);
      when "1001101111101" => q_unbuf <= my_rom(4989);
      when "1001101111110" => q_unbuf <= my_rom(4990);
      when "1001101111111" => q_unbuf <= my_rom(4991);
      when "1001110000000" => q_unbuf <= my_rom(4992);
      when "1001110000001" => q_unbuf <= my_rom(4993);
      when "1001110000010" => q_unbuf <= my_rom(4994);
      when "1001110000011" => q_unbuf <= my_rom(4995);
      when "1001110000100" => q_unbuf <= my_rom(4996);
      when "1001110000101" => q_unbuf <= my_rom(4997);
      when "1001110000110" => q_unbuf <= my_rom(4998);
      when "1001110000111" => q_unbuf <= my_rom(4999);
      when "1001110001000" => q_unbuf <= my_rom(5000);
      when "1001110001001" => q_unbuf <= my_rom(5001);
      when "1001110001010" => q_unbuf <= my_rom(5002);
      when "1001110001011" => q_unbuf <= my_rom(5003);
      when "1001110001100" => q_unbuf <= my_rom(5004);
      when "1001110001101" => q_unbuf <= my_rom(5005);
      when "1001110001110" => q_unbuf <= my_rom(5006);
      when "1001110001111" => q_unbuf <= my_rom(5007);
      when "1001110010000" => q_unbuf <= my_rom(5008);
      when "1001110010001" => q_unbuf <= my_rom(5009);
      when "1001110010010" => q_unbuf <= my_rom(5010);
      when "1001110010011" => q_unbuf <= my_rom(5011);
      when "1001110010100" => q_unbuf <= my_rom(5012);
      when "1001110010101" => q_unbuf <= my_rom(5013);
      when "1001110010110" => q_unbuf <= my_rom(5014);
      when "1001110010111" => q_unbuf <= my_rom(5015);
      when "1001110011000" => q_unbuf <= my_rom(5016);
      when "1001110011001" => q_unbuf <= my_rom(5017);
      when "1001110011010" => q_unbuf <= my_rom(5018);
      when "1001110011011" => q_unbuf <= my_rom(5019);
      when "1001110011100" => q_unbuf <= my_rom(5020);
      when "1001110011101" => q_unbuf <= my_rom(5021);
      when "1001110011110" => q_unbuf <= my_rom(5022);
      when "1001110011111" => q_unbuf <= my_rom(5023);
      when "1001110100000" => q_unbuf <= my_rom(5024);
      when "1001110100001" => q_unbuf <= my_rom(5025);
      when "1001110100010" => q_unbuf <= my_rom(5026);
      when "1001110100011" => q_unbuf <= my_rom(5027);
      when "1001110100100" => q_unbuf <= my_rom(5028);
      when "1001110100101" => q_unbuf <= my_rom(5029);
      when "1001110100110" => q_unbuf <= my_rom(5030);
      when "1001110100111" => q_unbuf <= my_rom(5031);
      when "1001110101000" => q_unbuf <= my_rom(5032);
      when "1001110101001" => q_unbuf <= my_rom(5033);
      when "1001110101010" => q_unbuf <= my_rom(5034);
      when "1001110101011" => q_unbuf <= my_rom(5035);
      when "1001110101100" => q_unbuf <= my_rom(5036);
      when "1001110101101" => q_unbuf <= my_rom(5037);
      when "1001110101110" => q_unbuf <= my_rom(5038);
      when "1001110101111" => q_unbuf <= my_rom(5039);
      when "1001110110000" => q_unbuf <= my_rom(5040);
      when "1001110110001" => q_unbuf <= my_rom(5041);
      when "1001110110010" => q_unbuf <= my_rom(5042);
      when "1001110110011" => q_unbuf <= my_rom(5043);
      when "1001110110100" => q_unbuf <= my_rom(5044);
      when "1001110110101" => q_unbuf <= my_rom(5045);
      when "1001110110110" => q_unbuf <= my_rom(5046);
      when "1001110110111" => q_unbuf <= my_rom(5047);
      when "1001110111000" => q_unbuf <= my_rom(5048);
      when "1001110111001" => q_unbuf <= my_rom(5049);
      when "1001110111010" => q_unbuf <= my_rom(5050);
      when "1001110111011" => q_unbuf <= my_rom(5051);
      when "1001110111100" => q_unbuf <= my_rom(5052);
      when "1001110111101" => q_unbuf <= my_rom(5053);
      when "1001110111110" => q_unbuf <= my_rom(5054);
      when "1001110111111" => q_unbuf <= my_rom(5055);
      when "1001111000000" => q_unbuf <= my_rom(5056);
      when "1001111000001" => q_unbuf <= my_rom(5057);
      when "1001111000010" => q_unbuf <= my_rom(5058);
      when "1001111000011" => q_unbuf <= my_rom(5059);
      when "1001111000100" => q_unbuf <= my_rom(5060);
      when "1001111000101" => q_unbuf <= my_rom(5061);
      when "1001111000110" => q_unbuf <= my_rom(5062);
      when "1001111000111" => q_unbuf <= my_rom(5063);
      when "1001111001000" => q_unbuf <= my_rom(5064);
      when "1001111001001" => q_unbuf <= my_rom(5065);
      when "1001111001010" => q_unbuf <= my_rom(5066);
      when "1001111001011" => q_unbuf <= my_rom(5067);
      when "1001111001100" => q_unbuf <= my_rom(5068);
      when "1001111001101" => q_unbuf <= my_rom(5069);
      when "1001111001110" => q_unbuf <= my_rom(5070);
      when "1001111001111" => q_unbuf <= my_rom(5071);
      when "1001111010000" => q_unbuf <= my_rom(5072);
      when "1001111010001" => q_unbuf <= my_rom(5073);
      when "1001111010010" => q_unbuf <= my_rom(5074);
      when "1001111010011" => q_unbuf <= my_rom(5075);
      when "1001111010100" => q_unbuf <= my_rom(5076);
      when "1001111010101" => q_unbuf <= my_rom(5077);
      when "1001111010110" => q_unbuf <= my_rom(5078);
      when "1001111010111" => q_unbuf <= my_rom(5079);
      when "1001111011000" => q_unbuf <= my_rom(5080);
      when "1001111011001" => q_unbuf <= my_rom(5081);
      when "1001111011010" => q_unbuf <= my_rom(5082);
      when "1001111011011" => q_unbuf <= my_rom(5083);
      when "1001111011100" => q_unbuf <= my_rom(5084);
      when "1001111011101" => q_unbuf <= my_rom(5085);
      when "1001111011110" => q_unbuf <= my_rom(5086);
      when "1001111011111" => q_unbuf <= my_rom(5087);
      when "1001111100000" => q_unbuf <= my_rom(5088);
      when "1001111100001" => q_unbuf <= my_rom(5089);
      when "1001111100010" => q_unbuf <= my_rom(5090);
      when "1001111100011" => q_unbuf <= my_rom(5091);
      when "1001111100100" => q_unbuf <= my_rom(5092);
      when "1001111100101" => q_unbuf <= my_rom(5093);
      when "1001111100110" => q_unbuf <= my_rom(5094);
      when "1001111100111" => q_unbuf <= my_rom(5095);
      when "1001111101000" => q_unbuf <= my_rom(5096);
      when "1001111101001" => q_unbuf <= my_rom(5097);
      when "1001111101010" => q_unbuf <= my_rom(5098);
      when "1001111101011" => q_unbuf <= my_rom(5099);
      when "1001111101100" => q_unbuf <= my_rom(5100);
      when "1001111101101" => q_unbuf <= my_rom(5101);
      when "1001111101110" => q_unbuf <= my_rom(5102);
      when "1001111101111" => q_unbuf <= my_rom(5103);
      when "1001111110000" => q_unbuf <= my_rom(5104);
      when "1001111110001" => q_unbuf <= my_rom(5105);
      when "1001111110010" => q_unbuf <= my_rom(5106);
      when "1001111110011" => q_unbuf <= my_rom(5107);
      when "1001111110100" => q_unbuf <= my_rom(5108);
      when "1001111110101" => q_unbuf <= my_rom(5109);
      when "1001111110110" => q_unbuf <= my_rom(5110);
      when "1001111110111" => q_unbuf <= my_rom(5111);
      when "1001111111000" => q_unbuf <= my_rom(5112);
      when "1001111111001" => q_unbuf <= my_rom(5113);
      when "1001111111010" => q_unbuf <= my_rom(5114);
      when "1001111111011" => q_unbuf <= my_rom(5115);
      when "1001111111100" => q_unbuf <= my_rom(5116);
      when "1001111111101" => q_unbuf <= my_rom(5117);
      when "1001111111110" => q_unbuf <= my_rom(5118);
      when "1001111111111" => q_unbuf <= my_rom(5119);
      when "1010000000000" => q_unbuf <= my_rom(5120);
      when "1010000000001" => q_unbuf <= my_rom(5121);
      when "1010000000010" => q_unbuf <= my_rom(5122);
      when "1010000000011" => q_unbuf <= my_rom(5123);
      when "1010000000100" => q_unbuf <= my_rom(5124);
      when "1010000000101" => q_unbuf <= my_rom(5125);
      when "1010000000110" => q_unbuf <= my_rom(5126);
      when "1010000000111" => q_unbuf <= my_rom(5127);
      when "1010000001000" => q_unbuf <= my_rom(5128);
      when "1010000001001" => q_unbuf <= my_rom(5129);
      when "1010000001010" => q_unbuf <= my_rom(5130);
      when "1010000001011" => q_unbuf <= my_rom(5131);
      when "1010000001100" => q_unbuf <= my_rom(5132);
      when "1010000001101" => q_unbuf <= my_rom(5133);
      when "1010000001110" => q_unbuf <= my_rom(5134);
      when "1010000001111" => q_unbuf <= my_rom(5135);
      when "1010000010000" => q_unbuf <= my_rom(5136);
      when "1010000010001" => q_unbuf <= my_rom(5137);
      when "1010000010010" => q_unbuf <= my_rom(5138);
      when "1010000010011" => q_unbuf <= my_rom(5139);
      when "1010000010100" => q_unbuf <= my_rom(5140);
      when "1010000010101" => q_unbuf <= my_rom(5141);
      when "1010000010110" => q_unbuf <= my_rom(5142);
      when "1010000010111" => q_unbuf <= my_rom(5143);
      when "1010000011000" => q_unbuf <= my_rom(5144);
      when "1010000011001" => q_unbuf <= my_rom(5145);
      when "1010000011010" => q_unbuf <= my_rom(5146);
      when "1010000011011" => q_unbuf <= my_rom(5147);
      when "1010000011100" => q_unbuf <= my_rom(5148);
      when "1010000011101" => q_unbuf <= my_rom(5149);
      when "1010000011110" => q_unbuf <= my_rom(5150);
      when "1010000011111" => q_unbuf <= my_rom(5151);
      when "1010000100000" => q_unbuf <= my_rom(5152);
      when "1010000100001" => q_unbuf <= my_rom(5153);
      when "1010000100010" => q_unbuf <= my_rom(5154);
      when "1010000100011" => q_unbuf <= my_rom(5155);
      when "1010000100100" => q_unbuf <= my_rom(5156);
      when "1010000100101" => q_unbuf <= my_rom(5157);
      when "1010000100110" => q_unbuf <= my_rom(5158);
      when "1010000100111" => q_unbuf <= my_rom(5159);
      when "1010000101000" => q_unbuf <= my_rom(5160);
      when "1010000101001" => q_unbuf <= my_rom(5161);
      when "1010000101010" => q_unbuf <= my_rom(5162);
      when "1010000101011" => q_unbuf <= my_rom(5163);
      when "1010000101100" => q_unbuf <= my_rom(5164);
      when "1010000101101" => q_unbuf <= my_rom(5165);
      when "1010000101110" => q_unbuf <= my_rom(5166);
      when "1010000101111" => q_unbuf <= my_rom(5167);
      when "1010000110000" => q_unbuf <= my_rom(5168);
      when "1010000110001" => q_unbuf <= my_rom(5169);
      when "1010000110010" => q_unbuf <= my_rom(5170);
      when "1010000110011" => q_unbuf <= my_rom(5171);
      when "1010000110100" => q_unbuf <= my_rom(5172);
      when "1010000110101" => q_unbuf <= my_rom(5173);
      when "1010000110110" => q_unbuf <= my_rom(5174);
      when "1010000110111" => q_unbuf <= my_rom(5175);
      when "1010000111000" => q_unbuf <= my_rom(5176);
      when "1010000111001" => q_unbuf <= my_rom(5177);
      when "1010000111010" => q_unbuf <= my_rom(5178);
      when "1010000111011" => q_unbuf <= my_rom(5179);
      when "1010000111100" => q_unbuf <= my_rom(5180);
      when "1010000111101" => q_unbuf <= my_rom(5181);
      when "1010000111110" => q_unbuf <= my_rom(5182);
      when "1010000111111" => q_unbuf <= my_rom(5183);
      when "1010001000000" => q_unbuf <= my_rom(5184);
      when "1010001000001" => q_unbuf <= my_rom(5185);
      when "1010001000010" => q_unbuf <= my_rom(5186);
      when "1010001000011" => q_unbuf <= my_rom(5187);
      when "1010001000100" => q_unbuf <= my_rom(5188);
      when "1010001000101" => q_unbuf <= my_rom(5189);
      when "1010001000110" => q_unbuf <= my_rom(5190);
      when "1010001000111" => q_unbuf <= my_rom(5191);
      when "1010001001000" => q_unbuf <= my_rom(5192);
      when "1010001001001" => q_unbuf <= my_rom(5193);
      when "1010001001010" => q_unbuf <= my_rom(5194);
      when "1010001001011" => q_unbuf <= my_rom(5195);
      when "1010001001100" => q_unbuf <= my_rom(5196);
      when "1010001001101" => q_unbuf <= my_rom(5197);
      when "1010001001110" => q_unbuf <= my_rom(5198);
      when "1010001001111" => q_unbuf <= my_rom(5199);
      when "1010001010000" => q_unbuf <= my_rom(5200);
      when "1010001010001" => q_unbuf <= my_rom(5201);
      when "1010001010010" => q_unbuf <= my_rom(5202);
      when "1010001010011" => q_unbuf <= my_rom(5203);
      when "1010001010100" => q_unbuf <= my_rom(5204);
      when "1010001010101" => q_unbuf <= my_rom(5205);
      when "1010001010110" => q_unbuf <= my_rom(5206);
      when "1010001010111" => q_unbuf <= my_rom(5207);
      when "1010001011000" => q_unbuf <= my_rom(5208);
      when "1010001011001" => q_unbuf <= my_rom(5209);
      when "1010001011010" => q_unbuf <= my_rom(5210);
      when "1010001011011" => q_unbuf <= my_rom(5211);
      when "1010001011100" => q_unbuf <= my_rom(5212);
      when "1010001011101" => q_unbuf <= my_rom(5213);
      when "1010001011110" => q_unbuf <= my_rom(5214);
      when "1010001011111" => q_unbuf <= my_rom(5215);
      when "1010001100000" => q_unbuf <= my_rom(5216);
      when "1010001100001" => q_unbuf <= my_rom(5217);
      when "1010001100010" => q_unbuf <= my_rom(5218);
      when "1010001100011" => q_unbuf <= my_rom(5219);
      when "1010001100100" => q_unbuf <= my_rom(5220);
      when "1010001100101" => q_unbuf <= my_rom(5221);
      when "1010001100110" => q_unbuf <= my_rom(5222);
      when "1010001100111" => q_unbuf <= my_rom(5223);
      when "1010001101000" => q_unbuf <= my_rom(5224);
      when "1010001101001" => q_unbuf <= my_rom(5225);
      when "1010001101010" => q_unbuf <= my_rom(5226);
      when "1010001101011" => q_unbuf <= my_rom(5227);
      when "1010001101100" => q_unbuf <= my_rom(5228);
      when "1010001101101" => q_unbuf <= my_rom(5229);
      when "1010001101110" => q_unbuf <= my_rom(5230);
      when "1010001101111" => q_unbuf <= my_rom(5231);
      when "1010001110000" => q_unbuf <= my_rom(5232);
      when "1010001110001" => q_unbuf <= my_rom(5233);
      when "1010001110010" => q_unbuf <= my_rom(5234);
      when "1010001110011" => q_unbuf <= my_rom(5235);
      when "1010001110100" => q_unbuf <= my_rom(5236);
      when "1010001110101" => q_unbuf <= my_rom(5237);
      when "1010001110110" => q_unbuf <= my_rom(5238);
      when "1010001110111" => q_unbuf <= my_rom(5239);
      when "1010001111000" => q_unbuf <= my_rom(5240);
      when "1010001111001" => q_unbuf <= my_rom(5241);
      when "1010001111010" => q_unbuf <= my_rom(5242);
      when "1010001111011" => q_unbuf <= my_rom(5243);
      when "1010001111100" => q_unbuf <= my_rom(5244);
      when "1010001111101" => q_unbuf <= my_rom(5245);
      when "1010001111110" => q_unbuf <= my_rom(5246);
      when "1010001111111" => q_unbuf <= my_rom(5247);
      when "1010010000000" => q_unbuf <= my_rom(5248);
      when "1010010000001" => q_unbuf <= my_rom(5249);
      when "1010010000010" => q_unbuf <= my_rom(5250);
      when "1010010000011" => q_unbuf <= my_rom(5251);
      when "1010010000100" => q_unbuf <= my_rom(5252);
      when "1010010000101" => q_unbuf <= my_rom(5253);
      when "1010010000110" => q_unbuf <= my_rom(5254);
      when "1010010000111" => q_unbuf <= my_rom(5255);
      when "1010010001000" => q_unbuf <= my_rom(5256);
      when "1010010001001" => q_unbuf <= my_rom(5257);
      when "1010010001010" => q_unbuf <= my_rom(5258);
      when "1010010001011" => q_unbuf <= my_rom(5259);
      when "1010010001100" => q_unbuf <= my_rom(5260);
      when "1010010001101" => q_unbuf <= my_rom(5261);
      when "1010010001110" => q_unbuf <= my_rom(5262);
      when "1010010001111" => q_unbuf <= my_rom(5263);
      when "1010010010000" => q_unbuf <= my_rom(5264);
      when "1010010010001" => q_unbuf <= my_rom(5265);
      when "1010010010010" => q_unbuf <= my_rom(5266);
      when "1010010010011" => q_unbuf <= my_rom(5267);
      when "1010010010100" => q_unbuf <= my_rom(5268);
      when "1010010010101" => q_unbuf <= my_rom(5269);
      when "1010010010110" => q_unbuf <= my_rom(5270);
      when "1010010010111" => q_unbuf <= my_rom(5271);
      when "1010010011000" => q_unbuf <= my_rom(5272);
      when "1010010011001" => q_unbuf <= my_rom(5273);
      when "1010010011010" => q_unbuf <= my_rom(5274);
      when "1010010011011" => q_unbuf <= my_rom(5275);
      when "1010010011100" => q_unbuf <= my_rom(5276);
      when "1010010011101" => q_unbuf <= my_rom(5277);
      when "1010010011110" => q_unbuf <= my_rom(5278);
      when "1010010011111" => q_unbuf <= my_rom(5279);
      when "1010010100000" => q_unbuf <= my_rom(5280);
      when "1010010100001" => q_unbuf <= my_rom(5281);
      when "1010010100010" => q_unbuf <= my_rom(5282);
      when "1010010100011" => q_unbuf <= my_rom(5283);
      when "1010010100100" => q_unbuf <= my_rom(5284);
      when "1010010100101" => q_unbuf <= my_rom(5285);
      when "1010010100110" => q_unbuf <= my_rom(5286);
      when "1010010100111" => q_unbuf <= my_rom(5287);
      when "1010010101000" => q_unbuf <= my_rom(5288);
      when "1010010101001" => q_unbuf <= my_rom(5289);
      when "1010010101010" => q_unbuf <= my_rom(5290);
      when "1010010101011" => q_unbuf <= my_rom(5291);
      when "1010010101100" => q_unbuf <= my_rom(5292);
      when "1010010101101" => q_unbuf <= my_rom(5293);
      when "1010010101110" => q_unbuf <= my_rom(5294);
      when "1010010101111" => q_unbuf <= my_rom(5295);
      when "1010010110000" => q_unbuf <= my_rom(5296);
      when "1010010110001" => q_unbuf <= my_rom(5297);
      when "1010010110010" => q_unbuf <= my_rom(5298);
      when "1010010110011" => q_unbuf <= my_rom(5299);
      when "1010010110100" => q_unbuf <= my_rom(5300);
      when "1010010110101" => q_unbuf <= my_rom(5301);
      when "1010010110110" => q_unbuf <= my_rom(5302);
      when "1010010110111" => q_unbuf <= my_rom(5303);
      when "1010010111000" => q_unbuf <= my_rom(5304);
      when "1010010111001" => q_unbuf <= my_rom(5305);
      when "1010010111010" => q_unbuf <= my_rom(5306);
      when "1010010111011" => q_unbuf <= my_rom(5307);
      when "1010010111100" => q_unbuf <= my_rom(5308);
      when "1010010111101" => q_unbuf <= my_rom(5309);
      when "1010010111110" => q_unbuf <= my_rom(5310);
      when "1010010111111" => q_unbuf <= my_rom(5311);
      when "1010011000000" => q_unbuf <= my_rom(5312);
      when "1010011000001" => q_unbuf <= my_rom(5313);
      when "1010011000010" => q_unbuf <= my_rom(5314);
      when "1010011000011" => q_unbuf <= my_rom(5315);
      when "1010011000100" => q_unbuf <= my_rom(5316);
      when "1010011000101" => q_unbuf <= my_rom(5317);
      when "1010011000110" => q_unbuf <= my_rom(5318);
      when "1010011000111" => q_unbuf <= my_rom(5319);
      when "1010011001000" => q_unbuf <= my_rom(5320);
      when "1010011001001" => q_unbuf <= my_rom(5321);
      when "1010011001010" => q_unbuf <= my_rom(5322);
      when "1010011001011" => q_unbuf <= my_rom(5323);
      when "1010011001100" => q_unbuf <= my_rom(5324);
      when "1010011001101" => q_unbuf <= my_rom(5325);
      when "1010011001110" => q_unbuf <= my_rom(5326);
      when "1010011001111" => q_unbuf <= my_rom(5327);
      when "1010011010000" => q_unbuf <= my_rom(5328);
      when "1010011010001" => q_unbuf <= my_rom(5329);
      when "1010011010010" => q_unbuf <= my_rom(5330);
      when "1010011010011" => q_unbuf <= my_rom(5331);
      when "1010011010100" => q_unbuf <= my_rom(5332);
      when "1010011010101" => q_unbuf <= my_rom(5333);
      when "1010011010110" => q_unbuf <= my_rom(5334);
      when "1010011010111" => q_unbuf <= my_rom(5335);
      when "1010011011000" => q_unbuf <= my_rom(5336);
      when "1010011011001" => q_unbuf <= my_rom(5337);
      when "1010011011010" => q_unbuf <= my_rom(5338);
      when "1010011011011" => q_unbuf <= my_rom(5339);
      when "1010011011100" => q_unbuf <= my_rom(5340);
      when "1010011011101" => q_unbuf <= my_rom(5341);
      when "1010011011110" => q_unbuf <= my_rom(5342);
      when "1010011011111" => q_unbuf <= my_rom(5343);
      when "1010011100000" => q_unbuf <= my_rom(5344);
      when "1010011100001" => q_unbuf <= my_rom(5345);
      when "1010011100010" => q_unbuf <= my_rom(5346);
      when "1010011100011" => q_unbuf <= my_rom(5347);
      when "1010011100100" => q_unbuf <= my_rom(5348);
      when "1010011100101" => q_unbuf <= my_rom(5349);
      when "1010011100110" => q_unbuf <= my_rom(5350);
      when "1010011100111" => q_unbuf <= my_rom(5351);
      when "1010011101000" => q_unbuf <= my_rom(5352);
      when "1010011101001" => q_unbuf <= my_rom(5353);
      when "1010011101010" => q_unbuf <= my_rom(5354);
      when "1010011101011" => q_unbuf <= my_rom(5355);
      when "1010011101100" => q_unbuf <= my_rom(5356);
      when "1010011101101" => q_unbuf <= my_rom(5357);
      when "1010011101110" => q_unbuf <= my_rom(5358);
      when "1010011101111" => q_unbuf <= my_rom(5359);
      when "1010011110000" => q_unbuf <= my_rom(5360);
      when "1010011110001" => q_unbuf <= my_rom(5361);
      when "1010011110010" => q_unbuf <= my_rom(5362);
      when "1010011110011" => q_unbuf <= my_rom(5363);
      when "1010011110100" => q_unbuf <= my_rom(5364);
      when "1010011110101" => q_unbuf <= my_rom(5365);
      when "1010011110110" => q_unbuf <= my_rom(5366);
      when "1010011110111" => q_unbuf <= my_rom(5367);
      when "1010011111000" => q_unbuf <= my_rom(5368);
      when "1010011111001" => q_unbuf <= my_rom(5369);
      when "1010011111010" => q_unbuf <= my_rom(5370);
      when "1010011111011" => q_unbuf <= my_rom(5371);
      when "1010011111100" => q_unbuf <= my_rom(5372);
      when "1010011111101" => q_unbuf <= my_rom(5373);
      when "1010011111110" => q_unbuf <= my_rom(5374);
      when "1010011111111" => q_unbuf <= my_rom(5375);
      when "1010100000000" => q_unbuf <= my_rom(5376);
      when "1010100000001" => q_unbuf <= my_rom(5377);
      when "1010100000010" => q_unbuf <= my_rom(5378);
      when "1010100000011" => q_unbuf <= my_rom(5379);
      when "1010100000100" => q_unbuf <= my_rom(5380);
      when "1010100000101" => q_unbuf <= my_rom(5381);
      when "1010100000110" => q_unbuf <= my_rom(5382);
      when "1010100000111" => q_unbuf <= my_rom(5383);
      when "1010100001000" => q_unbuf <= my_rom(5384);
      when "1010100001001" => q_unbuf <= my_rom(5385);
      when "1010100001010" => q_unbuf <= my_rom(5386);
      when "1010100001011" => q_unbuf <= my_rom(5387);
      when "1010100001100" => q_unbuf <= my_rom(5388);
      when "1010100001101" => q_unbuf <= my_rom(5389);
      when "1010100001110" => q_unbuf <= my_rom(5390);
      when "1010100001111" => q_unbuf <= my_rom(5391);
      when "1010100010000" => q_unbuf <= my_rom(5392);
      when "1010100010001" => q_unbuf <= my_rom(5393);
      when "1010100010010" => q_unbuf <= my_rom(5394);
      when "1010100010011" => q_unbuf <= my_rom(5395);
      when "1010100010100" => q_unbuf <= my_rom(5396);
      when "1010100010101" => q_unbuf <= my_rom(5397);
      when "1010100010110" => q_unbuf <= my_rom(5398);
      when "1010100010111" => q_unbuf <= my_rom(5399);
      when "1010100011000" => q_unbuf <= my_rom(5400);
      when "1010100011001" => q_unbuf <= my_rom(5401);
      when "1010100011010" => q_unbuf <= my_rom(5402);
      when "1010100011011" => q_unbuf <= my_rom(5403);
      when "1010100011100" => q_unbuf <= my_rom(5404);
      when "1010100011101" => q_unbuf <= my_rom(5405);
      when "1010100011110" => q_unbuf <= my_rom(5406);
      when "1010100011111" => q_unbuf <= my_rom(5407);
      when "1010100100000" => q_unbuf <= my_rom(5408);
      when "1010100100001" => q_unbuf <= my_rom(5409);
      when "1010100100010" => q_unbuf <= my_rom(5410);
      when "1010100100011" => q_unbuf <= my_rom(5411);
      when "1010100100100" => q_unbuf <= my_rom(5412);
      when "1010100100101" => q_unbuf <= my_rom(5413);
      when "1010100100110" => q_unbuf <= my_rom(5414);
      when "1010100100111" => q_unbuf <= my_rom(5415);
      when "1010100101000" => q_unbuf <= my_rom(5416);
      when "1010100101001" => q_unbuf <= my_rom(5417);
      when "1010100101010" => q_unbuf <= my_rom(5418);
      when "1010100101011" => q_unbuf <= my_rom(5419);
      when "1010100101100" => q_unbuf <= my_rom(5420);
      when "1010100101101" => q_unbuf <= my_rom(5421);
      when "1010100101110" => q_unbuf <= my_rom(5422);
      when "1010100101111" => q_unbuf <= my_rom(5423);
      when "1010100110000" => q_unbuf <= my_rom(5424);
      when "1010100110001" => q_unbuf <= my_rom(5425);
      when "1010100110010" => q_unbuf <= my_rom(5426);
      when "1010100110011" => q_unbuf <= my_rom(5427);
      when "1010100110100" => q_unbuf <= my_rom(5428);
      when "1010100110101" => q_unbuf <= my_rom(5429);
      when "1010100110110" => q_unbuf <= my_rom(5430);
      when "1010100110111" => q_unbuf <= my_rom(5431);
      when "1010100111000" => q_unbuf <= my_rom(5432);
      when "1010100111001" => q_unbuf <= my_rom(5433);
      when "1010100111010" => q_unbuf <= my_rom(5434);
      when "1010100111011" => q_unbuf <= my_rom(5435);
      when "1010100111100" => q_unbuf <= my_rom(5436);
      when "1010100111101" => q_unbuf <= my_rom(5437);
      when "1010100111110" => q_unbuf <= my_rom(5438);
      when "1010100111111" => q_unbuf <= my_rom(5439);
      when "1010101000000" => q_unbuf <= my_rom(5440);
      when "1010101000001" => q_unbuf <= my_rom(5441);
      when "1010101000010" => q_unbuf <= my_rom(5442);
      when "1010101000011" => q_unbuf <= my_rom(5443);
      when "1010101000100" => q_unbuf <= my_rom(5444);
      when "1010101000101" => q_unbuf <= my_rom(5445);
      when "1010101000110" => q_unbuf <= my_rom(5446);
      when "1010101000111" => q_unbuf <= my_rom(5447);
      when "1010101001000" => q_unbuf <= my_rom(5448);
      when "1010101001001" => q_unbuf <= my_rom(5449);
      when "1010101001010" => q_unbuf <= my_rom(5450);
      when "1010101001011" => q_unbuf <= my_rom(5451);
      when "1010101001100" => q_unbuf <= my_rom(5452);
      when "1010101001101" => q_unbuf <= my_rom(5453);
      when "1010101001110" => q_unbuf <= my_rom(5454);
      when "1010101001111" => q_unbuf <= my_rom(5455);
      when "1010101010000" => q_unbuf <= my_rom(5456);
      when "1010101010001" => q_unbuf <= my_rom(5457);
      when "1010101010010" => q_unbuf <= my_rom(5458);
      when "1010101010011" => q_unbuf <= my_rom(5459);
      when "1010101010100" => q_unbuf <= my_rom(5460);
      when "1010101010101" => q_unbuf <= my_rom(5461);
      when "1010101010110" => q_unbuf <= my_rom(5462);
      when "1010101010111" => q_unbuf <= my_rom(5463);
      when "1010101011000" => q_unbuf <= my_rom(5464);
      when "1010101011001" => q_unbuf <= my_rom(5465);
      when "1010101011010" => q_unbuf <= my_rom(5466);
      when "1010101011011" => q_unbuf <= my_rom(5467);
      when "1010101011100" => q_unbuf <= my_rom(5468);
      when "1010101011101" => q_unbuf <= my_rom(5469);
      when "1010101011110" => q_unbuf <= my_rom(5470);
      when "1010101011111" => q_unbuf <= my_rom(5471);
      when "1010101100000" => q_unbuf <= my_rom(5472);
      when "1010101100001" => q_unbuf <= my_rom(5473);
      when "1010101100010" => q_unbuf <= my_rom(5474);
      when "1010101100011" => q_unbuf <= my_rom(5475);
      when "1010101100100" => q_unbuf <= my_rom(5476);
      when "1010101100101" => q_unbuf <= my_rom(5477);
      when "1010101100110" => q_unbuf <= my_rom(5478);
      when "1010101100111" => q_unbuf <= my_rom(5479);
      when "1010101101000" => q_unbuf <= my_rom(5480);
      when "1010101101001" => q_unbuf <= my_rom(5481);
      when "1010101101010" => q_unbuf <= my_rom(5482);
      when "1010101101011" => q_unbuf <= my_rom(5483);
      when "1010101101100" => q_unbuf <= my_rom(5484);
      when "1010101101101" => q_unbuf <= my_rom(5485);
      when "1010101101110" => q_unbuf <= my_rom(5486);
      when "1010101101111" => q_unbuf <= my_rom(5487);
      when "1010101110000" => q_unbuf <= my_rom(5488);
      when "1010101110001" => q_unbuf <= my_rom(5489);
      when "1010101110010" => q_unbuf <= my_rom(5490);
      when "1010101110011" => q_unbuf <= my_rom(5491);
      when "1010101110100" => q_unbuf <= my_rom(5492);
      when "1010101110101" => q_unbuf <= my_rom(5493);
      when "1010101110110" => q_unbuf <= my_rom(5494);
      when "1010101110111" => q_unbuf <= my_rom(5495);
      when "1010101111000" => q_unbuf <= my_rom(5496);
      when "1010101111001" => q_unbuf <= my_rom(5497);
      when "1010101111010" => q_unbuf <= my_rom(5498);
      when "1010101111011" => q_unbuf <= my_rom(5499);
      when "1010101111100" => q_unbuf <= my_rom(5500);
      when "1010101111101" => q_unbuf <= my_rom(5501);
      when "1010101111110" => q_unbuf <= my_rom(5502);
      when "1010101111111" => q_unbuf <= my_rom(5503);
      when "1010110000000" => q_unbuf <= my_rom(5504);
      when "1010110000001" => q_unbuf <= my_rom(5505);
      when "1010110000010" => q_unbuf <= my_rom(5506);
      when "1010110000011" => q_unbuf <= my_rom(5507);
      when "1010110000100" => q_unbuf <= my_rom(5508);
      when "1010110000101" => q_unbuf <= my_rom(5509);
      when "1010110000110" => q_unbuf <= my_rom(5510);
      when "1010110000111" => q_unbuf <= my_rom(5511);
      when "1010110001000" => q_unbuf <= my_rom(5512);
      when "1010110001001" => q_unbuf <= my_rom(5513);
      when "1010110001010" => q_unbuf <= my_rom(5514);
      when "1010110001011" => q_unbuf <= my_rom(5515);
      when "1010110001100" => q_unbuf <= my_rom(5516);
      when "1010110001101" => q_unbuf <= my_rom(5517);
      when "1010110001110" => q_unbuf <= my_rom(5518);
      when "1010110001111" => q_unbuf <= my_rom(5519);
      when "1010110010000" => q_unbuf <= my_rom(5520);
      when "1010110010001" => q_unbuf <= my_rom(5521);
      when "1010110010010" => q_unbuf <= my_rom(5522);
      when "1010110010011" => q_unbuf <= my_rom(5523);
      when "1010110010100" => q_unbuf <= my_rom(5524);
      when "1010110010101" => q_unbuf <= my_rom(5525);
      when "1010110010110" => q_unbuf <= my_rom(5526);
      when "1010110010111" => q_unbuf <= my_rom(5527);
      when "1010110011000" => q_unbuf <= my_rom(5528);
      when "1010110011001" => q_unbuf <= my_rom(5529);
      when "1010110011010" => q_unbuf <= my_rom(5530);
      when "1010110011011" => q_unbuf <= my_rom(5531);
      when "1010110011100" => q_unbuf <= my_rom(5532);
      when "1010110011101" => q_unbuf <= my_rom(5533);
      when "1010110011110" => q_unbuf <= my_rom(5534);
      when "1010110011111" => q_unbuf <= my_rom(5535);
      when "1010110100000" => q_unbuf <= my_rom(5536);
      when "1010110100001" => q_unbuf <= my_rom(5537);
      when "1010110100010" => q_unbuf <= my_rom(5538);
      when "1010110100011" => q_unbuf <= my_rom(5539);
      when "1010110100100" => q_unbuf <= my_rom(5540);
      when "1010110100101" => q_unbuf <= my_rom(5541);
      when "1010110100110" => q_unbuf <= my_rom(5542);
      when "1010110100111" => q_unbuf <= my_rom(5543);
      when "1010110101000" => q_unbuf <= my_rom(5544);
      when "1010110101001" => q_unbuf <= my_rom(5545);
      when "1010110101010" => q_unbuf <= my_rom(5546);
      when "1010110101011" => q_unbuf <= my_rom(5547);
      when "1010110101100" => q_unbuf <= my_rom(5548);
      when "1010110101101" => q_unbuf <= my_rom(5549);
      when "1010110101110" => q_unbuf <= my_rom(5550);
      when "1010110101111" => q_unbuf <= my_rom(5551);
      when "1010110110000" => q_unbuf <= my_rom(5552);
      when "1010110110001" => q_unbuf <= my_rom(5553);
      when "1010110110010" => q_unbuf <= my_rom(5554);
      when "1010110110011" => q_unbuf <= my_rom(5555);
      when "1010110110100" => q_unbuf <= my_rom(5556);
      when "1010110110101" => q_unbuf <= my_rom(5557);
      when "1010110110110" => q_unbuf <= my_rom(5558);
      when "1010110110111" => q_unbuf <= my_rom(5559);
      when "1010110111000" => q_unbuf <= my_rom(5560);
      when "1010110111001" => q_unbuf <= my_rom(5561);
      when "1010110111010" => q_unbuf <= my_rom(5562);
      when "1010110111011" => q_unbuf <= my_rom(5563);
      when "1010110111100" => q_unbuf <= my_rom(5564);
      when "1010110111101" => q_unbuf <= my_rom(5565);
      when "1010110111110" => q_unbuf <= my_rom(5566);
      when "1010110111111" => q_unbuf <= my_rom(5567);
      when "1010111000000" => q_unbuf <= my_rom(5568);
      when "1010111000001" => q_unbuf <= my_rom(5569);
      when "1010111000010" => q_unbuf <= my_rom(5570);
      when "1010111000011" => q_unbuf <= my_rom(5571);
      when "1010111000100" => q_unbuf <= my_rom(5572);
      when "1010111000101" => q_unbuf <= my_rom(5573);
      when "1010111000110" => q_unbuf <= my_rom(5574);
      when "1010111000111" => q_unbuf <= my_rom(5575);
      when "1010111001000" => q_unbuf <= my_rom(5576);
      when "1010111001001" => q_unbuf <= my_rom(5577);
      when "1010111001010" => q_unbuf <= my_rom(5578);
      when "1010111001011" => q_unbuf <= my_rom(5579);
      when "1010111001100" => q_unbuf <= my_rom(5580);
      when "1010111001101" => q_unbuf <= my_rom(5581);
      when "1010111001110" => q_unbuf <= my_rom(5582);
      when "1010111001111" => q_unbuf <= my_rom(5583);
      when "1010111010000" => q_unbuf <= my_rom(5584);
      when "1010111010001" => q_unbuf <= my_rom(5585);
      when "1010111010010" => q_unbuf <= my_rom(5586);
      when "1010111010011" => q_unbuf <= my_rom(5587);
      when "1010111010100" => q_unbuf <= my_rom(5588);
      when "1010111010101" => q_unbuf <= my_rom(5589);
      when "1010111010110" => q_unbuf <= my_rom(5590);
      when "1010111010111" => q_unbuf <= my_rom(5591);
      when "1010111011000" => q_unbuf <= my_rom(5592);
      when "1010111011001" => q_unbuf <= my_rom(5593);
      when "1010111011010" => q_unbuf <= my_rom(5594);
      when "1010111011011" => q_unbuf <= my_rom(5595);
      when "1010111011100" => q_unbuf <= my_rom(5596);
      when "1010111011101" => q_unbuf <= my_rom(5597);
      when "1010111011110" => q_unbuf <= my_rom(5598);
      when "1010111011111" => q_unbuf <= my_rom(5599);
      when "1010111100000" => q_unbuf <= my_rom(5600);
      when "1010111100001" => q_unbuf <= my_rom(5601);
      when "1010111100010" => q_unbuf <= my_rom(5602);
      when "1010111100011" => q_unbuf <= my_rom(5603);
      when "1010111100100" => q_unbuf <= my_rom(5604);
      when "1010111100101" => q_unbuf <= my_rom(5605);
      when "1010111100110" => q_unbuf <= my_rom(5606);
      when "1010111100111" => q_unbuf <= my_rom(5607);
      when "1010111101000" => q_unbuf <= my_rom(5608);
      when "1010111101001" => q_unbuf <= my_rom(5609);
      when "1010111101010" => q_unbuf <= my_rom(5610);
      when "1010111101011" => q_unbuf <= my_rom(5611);
      when "1010111101100" => q_unbuf <= my_rom(5612);
      when "1010111101101" => q_unbuf <= my_rom(5613);
      when "1010111101110" => q_unbuf <= my_rom(5614);
      when "1010111101111" => q_unbuf <= my_rom(5615);
      when "1010111110000" => q_unbuf <= my_rom(5616);
      when "1010111110001" => q_unbuf <= my_rom(5617);
      when "1010111110010" => q_unbuf <= my_rom(5618);
      when "1010111110011" => q_unbuf <= my_rom(5619);
      when "1010111110100" => q_unbuf <= my_rom(5620);
      when "1010111110101" => q_unbuf <= my_rom(5621);
      when "1010111110110" => q_unbuf <= my_rom(5622);
      when "1010111110111" => q_unbuf <= my_rom(5623);
      when "1010111111000" => q_unbuf <= my_rom(5624);
      when "1010111111001" => q_unbuf <= my_rom(5625);
      when "1010111111010" => q_unbuf <= my_rom(5626);
      when "1010111111011" => q_unbuf <= my_rom(5627);
      when "1010111111100" => q_unbuf <= my_rom(5628);
      when "1010111111101" => q_unbuf <= my_rom(5629);
      when "1010111111110" => q_unbuf <= my_rom(5630);
      when "1010111111111" => q_unbuf <= my_rom(5631);
      when "1011000000000" => q_unbuf <= my_rom(5632);
      when "1011000000001" => q_unbuf <= my_rom(5633);
      when "1011000000010" => q_unbuf <= my_rom(5634);
      when "1011000000011" => q_unbuf <= my_rom(5635);
      when "1011000000100" => q_unbuf <= my_rom(5636);
      when "1011000000101" => q_unbuf <= my_rom(5637);
      when "1011000000110" => q_unbuf <= my_rom(5638);
      when "1011000000111" => q_unbuf <= my_rom(5639);
      when "1011000001000" => q_unbuf <= my_rom(5640);
      when "1011000001001" => q_unbuf <= my_rom(5641);
      when "1011000001010" => q_unbuf <= my_rom(5642);
      when "1011000001011" => q_unbuf <= my_rom(5643);
      when "1011000001100" => q_unbuf <= my_rom(5644);
      when "1011000001101" => q_unbuf <= my_rom(5645);
      when "1011000001110" => q_unbuf <= my_rom(5646);
      when "1011000001111" => q_unbuf <= my_rom(5647);
      when "1011000010000" => q_unbuf <= my_rom(5648);
      when "1011000010001" => q_unbuf <= my_rom(5649);
      when "1011000010010" => q_unbuf <= my_rom(5650);
      when "1011000010011" => q_unbuf <= my_rom(5651);
      when "1011000010100" => q_unbuf <= my_rom(5652);
      when "1011000010101" => q_unbuf <= my_rom(5653);
      when "1011000010110" => q_unbuf <= my_rom(5654);
      when "1011000010111" => q_unbuf <= my_rom(5655);
      when "1011000011000" => q_unbuf <= my_rom(5656);
      when "1011000011001" => q_unbuf <= my_rom(5657);
      when "1011000011010" => q_unbuf <= my_rom(5658);
      when "1011000011011" => q_unbuf <= my_rom(5659);
      when "1011000011100" => q_unbuf <= my_rom(5660);
      when "1011000011101" => q_unbuf <= my_rom(5661);
      when "1011000011110" => q_unbuf <= my_rom(5662);
      when "1011000011111" => q_unbuf <= my_rom(5663);
      when "1011000100000" => q_unbuf <= my_rom(5664);
      when "1011000100001" => q_unbuf <= my_rom(5665);
      when "1011000100010" => q_unbuf <= my_rom(5666);
      when "1011000100011" => q_unbuf <= my_rom(5667);
      when "1011000100100" => q_unbuf <= my_rom(5668);
      when "1011000100101" => q_unbuf <= my_rom(5669);
      when "1011000100110" => q_unbuf <= my_rom(5670);
      when "1011000100111" => q_unbuf <= my_rom(5671);
      when "1011000101000" => q_unbuf <= my_rom(5672);
      when "1011000101001" => q_unbuf <= my_rom(5673);
      when "1011000101010" => q_unbuf <= my_rom(5674);
      when "1011000101011" => q_unbuf <= my_rom(5675);
      when "1011000101100" => q_unbuf <= my_rom(5676);
      when "1011000101101" => q_unbuf <= my_rom(5677);
      when "1011000101110" => q_unbuf <= my_rom(5678);
      when "1011000101111" => q_unbuf <= my_rom(5679);
      when "1011000110000" => q_unbuf <= my_rom(5680);
      when "1011000110001" => q_unbuf <= my_rom(5681);
      when "1011000110010" => q_unbuf <= my_rom(5682);
      when "1011000110011" => q_unbuf <= my_rom(5683);
      when "1011000110100" => q_unbuf <= my_rom(5684);
      when "1011000110101" => q_unbuf <= my_rom(5685);
      when "1011000110110" => q_unbuf <= my_rom(5686);
      when "1011000110111" => q_unbuf <= my_rom(5687);
      when "1011000111000" => q_unbuf <= my_rom(5688);
      when "1011000111001" => q_unbuf <= my_rom(5689);
      when "1011000111010" => q_unbuf <= my_rom(5690);
      when "1011000111011" => q_unbuf <= my_rom(5691);
      when "1011000111100" => q_unbuf <= my_rom(5692);
      when "1011000111101" => q_unbuf <= my_rom(5693);
      when "1011000111110" => q_unbuf <= my_rom(5694);
      when "1011000111111" => q_unbuf <= my_rom(5695);
      when "1011001000000" => q_unbuf <= my_rom(5696);
      when "1011001000001" => q_unbuf <= my_rom(5697);
      when "1011001000010" => q_unbuf <= my_rom(5698);
      when "1011001000011" => q_unbuf <= my_rom(5699);
      when "1011001000100" => q_unbuf <= my_rom(5700);
      when "1011001000101" => q_unbuf <= my_rom(5701);
      when "1011001000110" => q_unbuf <= my_rom(5702);
      when "1011001000111" => q_unbuf <= my_rom(5703);
      when "1011001001000" => q_unbuf <= my_rom(5704);
      when "1011001001001" => q_unbuf <= my_rom(5705);
      when "1011001001010" => q_unbuf <= my_rom(5706);
      when "1011001001011" => q_unbuf <= my_rom(5707);
      when "1011001001100" => q_unbuf <= my_rom(5708);
      when "1011001001101" => q_unbuf <= my_rom(5709);
      when "1011001001110" => q_unbuf <= my_rom(5710);
      when "1011001001111" => q_unbuf <= my_rom(5711);
      when "1011001010000" => q_unbuf <= my_rom(5712);
      when "1011001010001" => q_unbuf <= my_rom(5713);
      when "1011001010010" => q_unbuf <= my_rom(5714);
      when "1011001010011" => q_unbuf <= my_rom(5715);
      when "1011001010100" => q_unbuf <= my_rom(5716);
      when "1011001010101" => q_unbuf <= my_rom(5717);
      when "1011001010110" => q_unbuf <= my_rom(5718);
      when "1011001010111" => q_unbuf <= my_rom(5719);
      when "1011001011000" => q_unbuf <= my_rom(5720);
      when "1011001011001" => q_unbuf <= my_rom(5721);
      when "1011001011010" => q_unbuf <= my_rom(5722);
      when "1011001011011" => q_unbuf <= my_rom(5723);
      when "1011001011100" => q_unbuf <= my_rom(5724);
      when "1011001011101" => q_unbuf <= my_rom(5725);
      when "1011001011110" => q_unbuf <= my_rom(5726);
      when "1011001011111" => q_unbuf <= my_rom(5727);
      when "1011001100000" => q_unbuf <= my_rom(5728);
      when "1011001100001" => q_unbuf <= my_rom(5729);
      when "1011001100010" => q_unbuf <= my_rom(5730);
      when "1011001100011" => q_unbuf <= my_rom(5731);
      when "1011001100100" => q_unbuf <= my_rom(5732);
      when "1011001100101" => q_unbuf <= my_rom(5733);
      when "1011001100110" => q_unbuf <= my_rom(5734);
      when "1011001100111" => q_unbuf <= my_rom(5735);
      when "1011001101000" => q_unbuf <= my_rom(5736);
      when "1011001101001" => q_unbuf <= my_rom(5737);
      when "1011001101010" => q_unbuf <= my_rom(5738);
      when "1011001101011" => q_unbuf <= my_rom(5739);
      when "1011001101100" => q_unbuf <= my_rom(5740);
      when "1011001101101" => q_unbuf <= my_rom(5741);
      when "1011001101110" => q_unbuf <= my_rom(5742);
      when "1011001101111" => q_unbuf <= my_rom(5743);
      when "1011001110000" => q_unbuf <= my_rom(5744);
      when "1011001110001" => q_unbuf <= my_rom(5745);
      when "1011001110010" => q_unbuf <= my_rom(5746);
      when "1011001110011" => q_unbuf <= my_rom(5747);
      when "1011001110100" => q_unbuf <= my_rom(5748);
      when "1011001110101" => q_unbuf <= my_rom(5749);
      when "1011001110110" => q_unbuf <= my_rom(5750);
      when "1011001110111" => q_unbuf <= my_rom(5751);
      when "1011001111000" => q_unbuf <= my_rom(5752);
      when "1011001111001" => q_unbuf <= my_rom(5753);
      when "1011001111010" => q_unbuf <= my_rom(5754);
      when "1011001111011" => q_unbuf <= my_rom(5755);
      when "1011001111100" => q_unbuf <= my_rom(5756);
      when "1011001111101" => q_unbuf <= my_rom(5757);
      when "1011001111110" => q_unbuf <= my_rom(5758);
      when "1011001111111" => q_unbuf <= my_rom(5759);
      when "1011010000000" => q_unbuf <= my_rom(5760);
      when "1011010000001" => q_unbuf <= my_rom(5761);
      when "1011010000010" => q_unbuf <= my_rom(5762);
      when "1011010000011" => q_unbuf <= my_rom(5763);
      when "1011010000100" => q_unbuf <= my_rom(5764);
      when "1011010000101" => q_unbuf <= my_rom(5765);
      when "1011010000110" => q_unbuf <= my_rom(5766);
      when "1011010000111" => q_unbuf <= my_rom(5767);
      when "1011010001000" => q_unbuf <= my_rom(5768);
      when "1011010001001" => q_unbuf <= my_rom(5769);
      when "1011010001010" => q_unbuf <= my_rom(5770);
      when "1011010001011" => q_unbuf <= my_rom(5771);
      when "1011010001100" => q_unbuf <= my_rom(5772);
      when "1011010001101" => q_unbuf <= my_rom(5773);
      when "1011010001110" => q_unbuf <= my_rom(5774);
      when "1011010001111" => q_unbuf <= my_rom(5775);
      when "1011010010000" => q_unbuf <= my_rom(5776);
      when "1011010010001" => q_unbuf <= my_rom(5777);
      when "1011010010010" => q_unbuf <= my_rom(5778);
      when "1011010010011" => q_unbuf <= my_rom(5779);
      when "1011010010100" => q_unbuf <= my_rom(5780);
      when "1011010010101" => q_unbuf <= my_rom(5781);
      when "1011010010110" => q_unbuf <= my_rom(5782);
      when "1011010010111" => q_unbuf <= my_rom(5783);
      when "1011010011000" => q_unbuf <= my_rom(5784);
      when "1011010011001" => q_unbuf <= my_rom(5785);
      when "1011010011010" => q_unbuf <= my_rom(5786);
      when "1011010011011" => q_unbuf <= my_rom(5787);
      when "1011010011100" => q_unbuf <= my_rom(5788);
      when "1011010011101" => q_unbuf <= my_rom(5789);
      when "1011010011110" => q_unbuf <= my_rom(5790);
      when "1011010011111" => q_unbuf <= my_rom(5791);
      when "1011010100000" => q_unbuf <= my_rom(5792);
      when "1011010100001" => q_unbuf <= my_rom(5793);
      when "1011010100010" => q_unbuf <= my_rom(5794);
      when "1011010100011" => q_unbuf <= my_rom(5795);
      when "1011010100100" => q_unbuf <= my_rom(5796);
      when "1011010100101" => q_unbuf <= my_rom(5797);
      when "1011010100110" => q_unbuf <= my_rom(5798);
      when "1011010100111" => q_unbuf <= my_rom(5799);
      when "1011010101000" => q_unbuf <= my_rom(5800);
      when "1011010101001" => q_unbuf <= my_rom(5801);
      when "1011010101010" => q_unbuf <= my_rom(5802);
      when "1011010101011" => q_unbuf <= my_rom(5803);
      when "1011010101100" => q_unbuf <= my_rom(5804);
      when "1011010101101" => q_unbuf <= my_rom(5805);
      when "1011010101110" => q_unbuf <= my_rom(5806);
      when "1011010101111" => q_unbuf <= my_rom(5807);
      when "1011010110000" => q_unbuf <= my_rom(5808);
      when "1011010110001" => q_unbuf <= my_rom(5809);
      when "1011010110010" => q_unbuf <= my_rom(5810);
      when "1011010110011" => q_unbuf <= my_rom(5811);
      when "1011010110100" => q_unbuf <= my_rom(5812);
      when "1011010110101" => q_unbuf <= my_rom(5813);
      when "1011010110110" => q_unbuf <= my_rom(5814);
      when "1011010110111" => q_unbuf <= my_rom(5815);
      when "1011010111000" => q_unbuf <= my_rom(5816);
      when "1011010111001" => q_unbuf <= my_rom(5817);
      when "1011010111010" => q_unbuf <= my_rom(5818);
      when "1011010111011" => q_unbuf <= my_rom(5819);
      when "1011010111100" => q_unbuf <= my_rom(5820);
      when "1011010111101" => q_unbuf <= my_rom(5821);
      when "1011010111110" => q_unbuf <= my_rom(5822);
      when "1011010111111" => q_unbuf <= my_rom(5823);
      when "1011011000000" => q_unbuf <= my_rom(5824);
      when "1011011000001" => q_unbuf <= my_rom(5825);
      when "1011011000010" => q_unbuf <= my_rom(5826);
      when "1011011000011" => q_unbuf <= my_rom(5827);
      when "1011011000100" => q_unbuf <= my_rom(5828);
      when "1011011000101" => q_unbuf <= my_rom(5829);
      when "1011011000110" => q_unbuf <= my_rom(5830);
      when "1011011000111" => q_unbuf <= my_rom(5831);
      when "1011011001000" => q_unbuf <= my_rom(5832);
      when "1011011001001" => q_unbuf <= my_rom(5833);
      when "1011011001010" => q_unbuf <= my_rom(5834);
      when "1011011001011" => q_unbuf <= my_rom(5835);
      when "1011011001100" => q_unbuf <= my_rom(5836);
      when "1011011001101" => q_unbuf <= my_rom(5837);
      when "1011011001110" => q_unbuf <= my_rom(5838);
      when "1011011001111" => q_unbuf <= my_rom(5839);
      when "1011011010000" => q_unbuf <= my_rom(5840);
      when "1011011010001" => q_unbuf <= my_rom(5841);
      when "1011011010010" => q_unbuf <= my_rom(5842);
      when "1011011010011" => q_unbuf <= my_rom(5843);
      when "1011011010100" => q_unbuf <= my_rom(5844);
      when "1011011010101" => q_unbuf <= my_rom(5845);
      when "1011011010110" => q_unbuf <= my_rom(5846);
      when "1011011010111" => q_unbuf <= my_rom(5847);
      when "1011011011000" => q_unbuf <= my_rom(5848);
      when "1011011011001" => q_unbuf <= my_rom(5849);
      when "1011011011010" => q_unbuf <= my_rom(5850);
      when "1011011011011" => q_unbuf <= my_rom(5851);
      when "1011011011100" => q_unbuf <= my_rom(5852);
      when "1011011011101" => q_unbuf <= my_rom(5853);
      when "1011011011110" => q_unbuf <= my_rom(5854);
      when "1011011011111" => q_unbuf <= my_rom(5855);
      when "1011011100000" => q_unbuf <= my_rom(5856);
      when "1011011100001" => q_unbuf <= my_rom(5857);
      when "1011011100010" => q_unbuf <= my_rom(5858);
      when "1011011100011" => q_unbuf <= my_rom(5859);
      when "1011011100100" => q_unbuf <= my_rom(5860);
      when "1011011100101" => q_unbuf <= my_rom(5861);
      when "1011011100110" => q_unbuf <= my_rom(5862);
      when "1011011100111" => q_unbuf <= my_rom(5863);
      when "1011011101000" => q_unbuf <= my_rom(5864);
      when "1011011101001" => q_unbuf <= my_rom(5865);
      when "1011011101010" => q_unbuf <= my_rom(5866);
      when "1011011101011" => q_unbuf <= my_rom(5867);
      when "1011011101100" => q_unbuf <= my_rom(5868);
      when "1011011101101" => q_unbuf <= my_rom(5869);
      when "1011011101110" => q_unbuf <= my_rom(5870);
      when "1011011101111" => q_unbuf <= my_rom(5871);
      when "1011011110000" => q_unbuf <= my_rom(5872);
      when "1011011110001" => q_unbuf <= my_rom(5873);
      when "1011011110010" => q_unbuf <= my_rom(5874);
      when "1011011110011" => q_unbuf <= my_rom(5875);
      when "1011011110100" => q_unbuf <= my_rom(5876);
      when "1011011110101" => q_unbuf <= my_rom(5877);
      when "1011011110110" => q_unbuf <= my_rom(5878);
      when "1011011110111" => q_unbuf <= my_rom(5879);
      when "1011011111000" => q_unbuf <= my_rom(5880);
      when "1011011111001" => q_unbuf <= my_rom(5881);
      when "1011011111010" => q_unbuf <= my_rom(5882);
      when "1011011111011" => q_unbuf <= my_rom(5883);
      when "1011011111100" => q_unbuf <= my_rom(5884);
      when "1011011111101" => q_unbuf <= my_rom(5885);
      when "1011011111110" => q_unbuf <= my_rom(5886);
      when "1011011111111" => q_unbuf <= my_rom(5887);
      when "1011100000000" => q_unbuf <= my_rom(5888);
      when "1011100000001" => q_unbuf <= my_rom(5889);
      when "1011100000010" => q_unbuf <= my_rom(5890);
      when "1011100000011" => q_unbuf <= my_rom(5891);
      when "1011100000100" => q_unbuf <= my_rom(5892);
      when "1011100000101" => q_unbuf <= my_rom(5893);
      when "1011100000110" => q_unbuf <= my_rom(5894);
      when "1011100000111" => q_unbuf <= my_rom(5895);
      when "1011100001000" => q_unbuf <= my_rom(5896);
      when "1011100001001" => q_unbuf <= my_rom(5897);
      when "1011100001010" => q_unbuf <= my_rom(5898);
      when "1011100001011" => q_unbuf <= my_rom(5899);
      when "1011100001100" => q_unbuf <= my_rom(5900);
      when "1011100001101" => q_unbuf <= my_rom(5901);
      when "1011100001110" => q_unbuf <= my_rom(5902);
      when "1011100001111" => q_unbuf <= my_rom(5903);
      when "1011100010000" => q_unbuf <= my_rom(5904);
      when "1011100010001" => q_unbuf <= my_rom(5905);
      when "1011100010010" => q_unbuf <= my_rom(5906);
      when "1011100010011" => q_unbuf <= my_rom(5907);
      when "1011100010100" => q_unbuf <= my_rom(5908);
      when "1011100010101" => q_unbuf <= my_rom(5909);
      when "1011100010110" => q_unbuf <= my_rom(5910);
      when "1011100010111" => q_unbuf <= my_rom(5911);
      when "1011100011000" => q_unbuf <= my_rom(5912);
      when "1011100011001" => q_unbuf <= my_rom(5913);
      when "1011100011010" => q_unbuf <= my_rom(5914);
      when "1011100011011" => q_unbuf <= my_rom(5915);
      when "1011100011100" => q_unbuf <= my_rom(5916);
      when "1011100011101" => q_unbuf <= my_rom(5917);
      when "1011100011110" => q_unbuf <= my_rom(5918);
      when "1011100011111" => q_unbuf <= my_rom(5919);
      when "1011100100000" => q_unbuf <= my_rom(5920);
      when "1011100100001" => q_unbuf <= my_rom(5921);
      when "1011100100010" => q_unbuf <= my_rom(5922);
      when "1011100100011" => q_unbuf <= my_rom(5923);
      when "1011100100100" => q_unbuf <= my_rom(5924);
      when "1011100100101" => q_unbuf <= my_rom(5925);
      when "1011100100110" => q_unbuf <= my_rom(5926);
      when "1011100100111" => q_unbuf <= my_rom(5927);
      when "1011100101000" => q_unbuf <= my_rom(5928);
      when "1011100101001" => q_unbuf <= my_rom(5929);
      when "1011100101010" => q_unbuf <= my_rom(5930);
      when "1011100101011" => q_unbuf <= my_rom(5931);
      when "1011100101100" => q_unbuf <= my_rom(5932);
      when "1011100101101" => q_unbuf <= my_rom(5933);
      when "1011100101110" => q_unbuf <= my_rom(5934);
      when "1011100101111" => q_unbuf <= my_rom(5935);
      when "1011100110000" => q_unbuf <= my_rom(5936);
      when "1011100110001" => q_unbuf <= my_rom(5937);
      when "1011100110010" => q_unbuf <= my_rom(5938);
      when "1011100110011" => q_unbuf <= my_rom(5939);
      when "1011100110100" => q_unbuf <= my_rom(5940);
      when "1011100110101" => q_unbuf <= my_rom(5941);
      when "1011100110110" => q_unbuf <= my_rom(5942);
      when "1011100110111" => q_unbuf <= my_rom(5943);
      when "1011100111000" => q_unbuf <= my_rom(5944);
      when "1011100111001" => q_unbuf <= my_rom(5945);
      when "1011100111010" => q_unbuf <= my_rom(5946);
      when "1011100111011" => q_unbuf <= my_rom(5947);
      when "1011100111100" => q_unbuf <= my_rom(5948);
      when "1011100111101" => q_unbuf <= my_rom(5949);
      when "1011100111110" => q_unbuf <= my_rom(5950);
      when "1011100111111" => q_unbuf <= my_rom(5951);
      when "1011101000000" => q_unbuf <= my_rom(5952);
      when "1011101000001" => q_unbuf <= my_rom(5953);
      when "1011101000010" => q_unbuf <= my_rom(5954);
      when "1011101000011" => q_unbuf <= my_rom(5955);
      when "1011101000100" => q_unbuf <= my_rom(5956);
      when "1011101000101" => q_unbuf <= my_rom(5957);
      when "1011101000110" => q_unbuf <= my_rom(5958);
      when "1011101000111" => q_unbuf <= my_rom(5959);
      when "1011101001000" => q_unbuf <= my_rom(5960);
      when "1011101001001" => q_unbuf <= my_rom(5961);
      when "1011101001010" => q_unbuf <= my_rom(5962);
      when "1011101001011" => q_unbuf <= my_rom(5963);
      when "1011101001100" => q_unbuf <= my_rom(5964);
      when "1011101001101" => q_unbuf <= my_rom(5965);
      when "1011101001110" => q_unbuf <= my_rom(5966);
      when "1011101001111" => q_unbuf <= my_rom(5967);
      when "1011101010000" => q_unbuf <= my_rom(5968);
      when "1011101010001" => q_unbuf <= my_rom(5969);
      when "1011101010010" => q_unbuf <= my_rom(5970);
      when "1011101010011" => q_unbuf <= my_rom(5971);
      when "1011101010100" => q_unbuf <= my_rom(5972);
      when "1011101010101" => q_unbuf <= my_rom(5973);
      when "1011101010110" => q_unbuf <= my_rom(5974);
      when "1011101010111" => q_unbuf <= my_rom(5975);
      when "1011101011000" => q_unbuf <= my_rom(5976);
      when "1011101011001" => q_unbuf <= my_rom(5977);
      when "1011101011010" => q_unbuf <= my_rom(5978);
      when "1011101011011" => q_unbuf <= my_rom(5979);
      when "1011101011100" => q_unbuf <= my_rom(5980);
      when "1011101011101" => q_unbuf <= my_rom(5981);
      when "1011101011110" => q_unbuf <= my_rom(5982);
      when "1011101011111" => q_unbuf <= my_rom(5983);
      when "1011101100000" => q_unbuf <= my_rom(5984);
      when "1011101100001" => q_unbuf <= my_rom(5985);
      when "1011101100010" => q_unbuf <= my_rom(5986);
      when "1011101100011" => q_unbuf <= my_rom(5987);
      when "1011101100100" => q_unbuf <= my_rom(5988);
      when "1011101100101" => q_unbuf <= my_rom(5989);
      when "1011101100110" => q_unbuf <= my_rom(5990);
      when "1011101100111" => q_unbuf <= my_rom(5991);
      when "1011101101000" => q_unbuf <= my_rom(5992);
      when "1011101101001" => q_unbuf <= my_rom(5993);
      when "1011101101010" => q_unbuf <= my_rom(5994);
      when "1011101101011" => q_unbuf <= my_rom(5995);
      when "1011101101100" => q_unbuf <= my_rom(5996);
      when "1011101101101" => q_unbuf <= my_rom(5997);
      when "1011101101110" => q_unbuf <= my_rom(5998);
      when "1011101101111" => q_unbuf <= my_rom(5999);
      when "1011101110000" => q_unbuf <= my_rom(6000);
      when "1011101110001" => q_unbuf <= my_rom(6001);
      when "1011101110010" => q_unbuf <= my_rom(6002);
      when "1011101110011" => q_unbuf <= my_rom(6003);
      when "1011101110100" => q_unbuf <= my_rom(6004);
      when "1011101110101" => q_unbuf <= my_rom(6005);
      when "1011101110110" => q_unbuf <= my_rom(6006);
      when "1011101110111" => q_unbuf <= my_rom(6007);
      when "1011101111000" => q_unbuf <= my_rom(6008);
      when "1011101111001" => q_unbuf <= my_rom(6009);
      when "1011101111010" => q_unbuf <= my_rom(6010);
      when "1011101111011" => q_unbuf <= my_rom(6011);
      when "1011101111100" => q_unbuf <= my_rom(6012);
      when "1011101111101" => q_unbuf <= my_rom(6013);
      when "1011101111110" => q_unbuf <= my_rom(6014);
      when "1011101111111" => q_unbuf <= my_rom(6015);
      when "1011110000000" => q_unbuf <= my_rom(6016);
      when "1011110000001" => q_unbuf <= my_rom(6017);
      when "1011110000010" => q_unbuf <= my_rom(6018);
      when "1011110000011" => q_unbuf <= my_rom(6019);
      when "1011110000100" => q_unbuf <= my_rom(6020);
      when "1011110000101" => q_unbuf <= my_rom(6021);
      when "1011110000110" => q_unbuf <= my_rom(6022);
      when "1011110000111" => q_unbuf <= my_rom(6023);
      when "1011110001000" => q_unbuf <= my_rom(6024);
      when "1011110001001" => q_unbuf <= my_rom(6025);
      when "1011110001010" => q_unbuf <= my_rom(6026);
      when "1011110001011" => q_unbuf <= my_rom(6027);
      when "1011110001100" => q_unbuf <= my_rom(6028);
      when "1011110001101" => q_unbuf <= my_rom(6029);
      when "1011110001110" => q_unbuf <= my_rom(6030);
      when "1011110001111" => q_unbuf <= my_rom(6031);
      when "1011110010000" => q_unbuf <= my_rom(6032);
      when "1011110010001" => q_unbuf <= my_rom(6033);
      when "1011110010010" => q_unbuf <= my_rom(6034);
      when "1011110010011" => q_unbuf <= my_rom(6035);
      when "1011110010100" => q_unbuf <= my_rom(6036);
      when "1011110010101" => q_unbuf <= my_rom(6037);
      when "1011110010110" => q_unbuf <= my_rom(6038);
      when "1011110010111" => q_unbuf <= my_rom(6039);
      when "1011110011000" => q_unbuf <= my_rom(6040);
      when "1011110011001" => q_unbuf <= my_rom(6041);
      when "1011110011010" => q_unbuf <= my_rom(6042);
      when "1011110011011" => q_unbuf <= my_rom(6043);
      when "1011110011100" => q_unbuf <= my_rom(6044);
      when "1011110011101" => q_unbuf <= my_rom(6045);
      when "1011110011110" => q_unbuf <= my_rom(6046);
      when "1011110011111" => q_unbuf <= my_rom(6047);
      when "1011110100000" => q_unbuf <= my_rom(6048);
      when "1011110100001" => q_unbuf <= my_rom(6049);
      when "1011110100010" => q_unbuf <= my_rom(6050);
      when "1011110100011" => q_unbuf <= my_rom(6051);
      when "1011110100100" => q_unbuf <= my_rom(6052);
      when "1011110100101" => q_unbuf <= my_rom(6053);
      when "1011110100110" => q_unbuf <= my_rom(6054);
      when "1011110100111" => q_unbuf <= my_rom(6055);
      when "1011110101000" => q_unbuf <= my_rom(6056);
      when "1011110101001" => q_unbuf <= my_rom(6057);
      when "1011110101010" => q_unbuf <= my_rom(6058);
      when "1011110101011" => q_unbuf <= my_rom(6059);
      when "1011110101100" => q_unbuf <= my_rom(6060);
      when "1011110101101" => q_unbuf <= my_rom(6061);
      when "1011110101110" => q_unbuf <= my_rom(6062);
      when "1011110101111" => q_unbuf <= my_rom(6063);
      when "1011110110000" => q_unbuf <= my_rom(6064);
      when "1011110110001" => q_unbuf <= my_rom(6065);
      when "1011110110010" => q_unbuf <= my_rom(6066);
      when "1011110110011" => q_unbuf <= my_rom(6067);
      when "1011110110100" => q_unbuf <= my_rom(6068);
      when "1011110110101" => q_unbuf <= my_rom(6069);
      when "1011110110110" => q_unbuf <= my_rom(6070);
      when "1011110110111" => q_unbuf <= my_rom(6071);
      when "1011110111000" => q_unbuf <= my_rom(6072);
      when "1011110111001" => q_unbuf <= my_rom(6073);
      when "1011110111010" => q_unbuf <= my_rom(6074);
      when "1011110111011" => q_unbuf <= my_rom(6075);
      when "1011110111100" => q_unbuf <= my_rom(6076);
      when "1011110111101" => q_unbuf <= my_rom(6077);
      when "1011110111110" => q_unbuf <= my_rom(6078);
      when "1011110111111" => q_unbuf <= my_rom(6079);
      when "1011111000000" => q_unbuf <= my_rom(6080);
      when "1011111000001" => q_unbuf <= my_rom(6081);
      when "1011111000010" => q_unbuf <= my_rom(6082);
      when "1011111000011" => q_unbuf <= my_rom(6083);
      when "1011111000100" => q_unbuf <= my_rom(6084);
      when "1011111000101" => q_unbuf <= my_rom(6085);
      when "1011111000110" => q_unbuf <= my_rom(6086);
      when "1011111000111" => q_unbuf <= my_rom(6087);
      when "1011111001000" => q_unbuf <= my_rom(6088);
      when "1011111001001" => q_unbuf <= my_rom(6089);
      when "1011111001010" => q_unbuf <= my_rom(6090);
      when "1011111001011" => q_unbuf <= my_rom(6091);
      when "1011111001100" => q_unbuf <= my_rom(6092);
      when "1011111001101" => q_unbuf <= my_rom(6093);
      when "1011111001110" => q_unbuf <= my_rom(6094);
      when "1011111001111" => q_unbuf <= my_rom(6095);
      when "1011111010000" => q_unbuf <= my_rom(6096);
      when "1011111010001" => q_unbuf <= my_rom(6097);
      when "1011111010010" => q_unbuf <= my_rom(6098);
      when "1011111010011" => q_unbuf <= my_rom(6099);
      when "1011111010100" => q_unbuf <= my_rom(6100);
      when "1011111010101" => q_unbuf <= my_rom(6101);
      when "1011111010110" => q_unbuf <= my_rom(6102);
      when "1011111010111" => q_unbuf <= my_rom(6103);
      when "1011111011000" => q_unbuf <= my_rom(6104);
      when "1011111011001" => q_unbuf <= my_rom(6105);
      when "1011111011010" => q_unbuf <= my_rom(6106);
      when "1011111011011" => q_unbuf <= my_rom(6107);
      when "1011111011100" => q_unbuf <= my_rom(6108);
      when "1011111011101" => q_unbuf <= my_rom(6109);
      when "1011111011110" => q_unbuf <= my_rom(6110);
      when "1011111011111" => q_unbuf <= my_rom(6111);
      when "1011111100000" => q_unbuf <= my_rom(6112);
      when "1011111100001" => q_unbuf <= my_rom(6113);
      when "1011111100010" => q_unbuf <= my_rom(6114);
      when "1011111100011" => q_unbuf <= my_rom(6115);
      when "1011111100100" => q_unbuf <= my_rom(6116);
      when "1011111100101" => q_unbuf <= my_rom(6117);
      when "1011111100110" => q_unbuf <= my_rom(6118);
      when "1011111100111" => q_unbuf <= my_rom(6119);
      when "1011111101000" => q_unbuf <= my_rom(6120);
      when "1011111101001" => q_unbuf <= my_rom(6121);
      when "1011111101010" => q_unbuf <= my_rom(6122);
      when "1011111101011" => q_unbuf <= my_rom(6123);
      when "1011111101100" => q_unbuf <= my_rom(6124);
      when "1011111101101" => q_unbuf <= my_rom(6125);
      when "1011111101110" => q_unbuf <= my_rom(6126);
      when "1011111101111" => q_unbuf <= my_rom(6127);
      when "1011111110000" => q_unbuf <= my_rom(6128);
      when "1011111110001" => q_unbuf <= my_rom(6129);
      when "1011111110010" => q_unbuf <= my_rom(6130);
      when "1011111110011" => q_unbuf <= my_rom(6131);
      when "1011111110100" => q_unbuf <= my_rom(6132);
      when "1011111110101" => q_unbuf <= my_rom(6133);
      when "1011111110110" => q_unbuf <= my_rom(6134);
      when "1011111110111" => q_unbuf <= my_rom(6135);
      when "1011111111000" => q_unbuf <= my_rom(6136);
      when "1011111111001" => q_unbuf <= my_rom(6137);
      when "1011111111010" => q_unbuf <= my_rom(6138);
      when "1011111111011" => q_unbuf <= my_rom(6139);
      when "1011111111100" => q_unbuf <= my_rom(6140);
      when "1011111111101" => q_unbuf <= my_rom(6141);
      when "1011111111110" => q_unbuf <= my_rom(6142);
      when "1011111111111" => q_unbuf <= my_rom(6143);
      when "1100000000000" => q_unbuf <= my_rom(6144);
      when "1100000000001" => q_unbuf <= my_rom(6145);
      when "1100000000010" => q_unbuf <= my_rom(6146);
      when "1100000000011" => q_unbuf <= my_rom(6147);
      when "1100000000100" => q_unbuf <= my_rom(6148);
      when "1100000000101" => q_unbuf <= my_rom(6149);
      when "1100000000110" => q_unbuf <= my_rom(6150);
      when "1100000000111" => q_unbuf <= my_rom(6151);
      when "1100000001000" => q_unbuf <= my_rom(6152);
      when "1100000001001" => q_unbuf <= my_rom(6153);
      when "1100000001010" => q_unbuf <= my_rom(6154);
      when "1100000001011" => q_unbuf <= my_rom(6155);
      when "1100000001100" => q_unbuf <= my_rom(6156);
      when "1100000001101" => q_unbuf <= my_rom(6157);
      when "1100000001110" => q_unbuf <= my_rom(6158);
      when "1100000001111" => q_unbuf <= my_rom(6159);
      when "1100000010000" => q_unbuf <= my_rom(6160);
      when "1100000010001" => q_unbuf <= my_rom(6161);
      when "1100000010010" => q_unbuf <= my_rom(6162);
      when "1100000010011" => q_unbuf <= my_rom(6163);
      when "1100000010100" => q_unbuf <= my_rom(6164);
      when "1100000010101" => q_unbuf <= my_rom(6165);
      when "1100000010110" => q_unbuf <= my_rom(6166);
      when "1100000010111" => q_unbuf <= my_rom(6167);
      when "1100000011000" => q_unbuf <= my_rom(6168);
      when "1100000011001" => q_unbuf <= my_rom(6169);
      when "1100000011010" => q_unbuf <= my_rom(6170);
      when "1100000011011" => q_unbuf <= my_rom(6171);
      when "1100000011100" => q_unbuf <= my_rom(6172);
      when "1100000011101" => q_unbuf <= my_rom(6173);
      when "1100000011110" => q_unbuf <= my_rom(6174);
      when "1100000011111" => q_unbuf <= my_rom(6175);
      when "1100000100000" => q_unbuf <= my_rom(6176);
      when "1100000100001" => q_unbuf <= my_rom(6177);
      when "1100000100010" => q_unbuf <= my_rom(6178);
      when "1100000100011" => q_unbuf <= my_rom(6179);
      when "1100000100100" => q_unbuf <= my_rom(6180);
      when "1100000100101" => q_unbuf <= my_rom(6181);
      when "1100000100110" => q_unbuf <= my_rom(6182);
      when "1100000100111" => q_unbuf <= my_rom(6183);
      when "1100000101000" => q_unbuf <= my_rom(6184);
      when "1100000101001" => q_unbuf <= my_rom(6185);
      when "1100000101010" => q_unbuf <= my_rom(6186);
      when "1100000101011" => q_unbuf <= my_rom(6187);
      when "1100000101100" => q_unbuf <= my_rom(6188);
      when "1100000101101" => q_unbuf <= my_rom(6189);
      when "1100000101110" => q_unbuf <= my_rom(6190);
      when "1100000101111" => q_unbuf <= my_rom(6191);
      when "1100000110000" => q_unbuf <= my_rom(6192);
      when "1100000110001" => q_unbuf <= my_rom(6193);
      when "1100000110010" => q_unbuf <= my_rom(6194);
      when "1100000110011" => q_unbuf <= my_rom(6195);
      when "1100000110100" => q_unbuf <= my_rom(6196);
      when "1100000110101" => q_unbuf <= my_rom(6197);
      when "1100000110110" => q_unbuf <= my_rom(6198);
      when "1100000110111" => q_unbuf <= my_rom(6199);
      when "1100000111000" => q_unbuf <= my_rom(6200);
      when "1100000111001" => q_unbuf <= my_rom(6201);
      when "1100000111010" => q_unbuf <= my_rom(6202);
      when "1100000111011" => q_unbuf <= my_rom(6203);
      when "1100000111100" => q_unbuf <= my_rom(6204);
      when "1100000111101" => q_unbuf <= my_rom(6205);
      when "1100000111110" => q_unbuf <= my_rom(6206);
      when "1100000111111" => q_unbuf <= my_rom(6207);
      when "1100001000000" => q_unbuf <= my_rom(6208);
      when "1100001000001" => q_unbuf <= my_rom(6209);
      when "1100001000010" => q_unbuf <= my_rom(6210);
      when "1100001000011" => q_unbuf <= my_rom(6211);
      when "1100001000100" => q_unbuf <= my_rom(6212);
      when "1100001000101" => q_unbuf <= my_rom(6213);
      when "1100001000110" => q_unbuf <= my_rom(6214);
      when "1100001000111" => q_unbuf <= my_rom(6215);
      when "1100001001000" => q_unbuf <= my_rom(6216);
      when "1100001001001" => q_unbuf <= my_rom(6217);
      when "1100001001010" => q_unbuf <= my_rom(6218);
      when "1100001001011" => q_unbuf <= my_rom(6219);
      when "1100001001100" => q_unbuf <= my_rom(6220);
      when "1100001001101" => q_unbuf <= my_rom(6221);
      when "1100001001110" => q_unbuf <= my_rom(6222);
      when "1100001001111" => q_unbuf <= my_rom(6223);
      when "1100001010000" => q_unbuf <= my_rom(6224);
      when "1100001010001" => q_unbuf <= my_rom(6225);
      when "1100001010010" => q_unbuf <= my_rom(6226);
      when "1100001010011" => q_unbuf <= my_rom(6227);
      when "1100001010100" => q_unbuf <= my_rom(6228);
      when "1100001010101" => q_unbuf <= my_rom(6229);
      when "1100001010110" => q_unbuf <= my_rom(6230);
      when "1100001010111" => q_unbuf <= my_rom(6231);
      when "1100001011000" => q_unbuf <= my_rom(6232);
      when "1100001011001" => q_unbuf <= my_rom(6233);
      when "1100001011010" => q_unbuf <= my_rom(6234);
      when "1100001011011" => q_unbuf <= my_rom(6235);
      when "1100001011100" => q_unbuf <= my_rom(6236);
      when "1100001011101" => q_unbuf <= my_rom(6237);
      when "1100001011110" => q_unbuf <= my_rom(6238);
      when "1100001011111" => q_unbuf <= my_rom(6239);
      when "1100001100000" => q_unbuf <= my_rom(6240);
      when "1100001100001" => q_unbuf <= my_rom(6241);
      when "1100001100010" => q_unbuf <= my_rom(6242);
      when "1100001100011" => q_unbuf <= my_rom(6243);
      when "1100001100100" => q_unbuf <= my_rom(6244);
      when "1100001100101" => q_unbuf <= my_rom(6245);
      when "1100001100110" => q_unbuf <= my_rom(6246);
      when "1100001100111" => q_unbuf <= my_rom(6247);
      when "1100001101000" => q_unbuf <= my_rom(6248);
      when "1100001101001" => q_unbuf <= my_rom(6249);
      when "1100001101010" => q_unbuf <= my_rom(6250);
      when "1100001101011" => q_unbuf <= my_rom(6251);
      when "1100001101100" => q_unbuf <= my_rom(6252);
      when "1100001101101" => q_unbuf <= my_rom(6253);
      when "1100001101110" => q_unbuf <= my_rom(6254);
      when "1100001101111" => q_unbuf <= my_rom(6255);
      when "1100001110000" => q_unbuf <= my_rom(6256);
      when "1100001110001" => q_unbuf <= my_rom(6257);
      when "1100001110010" => q_unbuf <= my_rom(6258);
      when "1100001110011" => q_unbuf <= my_rom(6259);
      when "1100001110100" => q_unbuf <= my_rom(6260);
      when "1100001110101" => q_unbuf <= my_rom(6261);
      when "1100001110110" => q_unbuf <= my_rom(6262);
      when "1100001110111" => q_unbuf <= my_rom(6263);
      when "1100001111000" => q_unbuf <= my_rom(6264);
      when "1100001111001" => q_unbuf <= my_rom(6265);
      when "1100001111010" => q_unbuf <= my_rom(6266);
      when "1100001111011" => q_unbuf <= my_rom(6267);
      when "1100001111100" => q_unbuf <= my_rom(6268);
      when "1100001111101" => q_unbuf <= my_rom(6269);
      when "1100001111110" => q_unbuf <= my_rom(6270);
      when "1100001111111" => q_unbuf <= my_rom(6271);
      when "1100010000000" => q_unbuf <= my_rom(6272);
      when "1100010000001" => q_unbuf <= my_rom(6273);
      when "1100010000010" => q_unbuf <= my_rom(6274);
      when "1100010000011" => q_unbuf <= my_rom(6275);
      when "1100010000100" => q_unbuf <= my_rom(6276);
      when "1100010000101" => q_unbuf <= my_rom(6277);
      when "1100010000110" => q_unbuf <= my_rom(6278);
      when "1100010000111" => q_unbuf <= my_rom(6279);
      when "1100010001000" => q_unbuf <= my_rom(6280);
      when "1100010001001" => q_unbuf <= my_rom(6281);
      when "1100010001010" => q_unbuf <= my_rom(6282);
      when "1100010001011" => q_unbuf <= my_rom(6283);
      when "1100010001100" => q_unbuf <= my_rom(6284);
      when "1100010001101" => q_unbuf <= my_rom(6285);
      when "1100010001110" => q_unbuf <= my_rom(6286);
      when "1100010001111" => q_unbuf <= my_rom(6287);
      when "1100010010000" => q_unbuf <= my_rom(6288);
      when "1100010010001" => q_unbuf <= my_rom(6289);
      when "1100010010010" => q_unbuf <= my_rom(6290);
      when "1100010010011" => q_unbuf <= my_rom(6291);
      when "1100010010100" => q_unbuf <= my_rom(6292);
      when "1100010010101" => q_unbuf <= my_rom(6293);
      when "1100010010110" => q_unbuf <= my_rom(6294);
      when "1100010010111" => q_unbuf <= my_rom(6295);
      when "1100010011000" => q_unbuf <= my_rom(6296);
      when "1100010011001" => q_unbuf <= my_rom(6297);
      when "1100010011010" => q_unbuf <= my_rom(6298);
      when "1100010011011" => q_unbuf <= my_rom(6299);
      when "1100010011100" => q_unbuf <= my_rom(6300);
      when "1100010011101" => q_unbuf <= my_rom(6301);
      when "1100010011110" => q_unbuf <= my_rom(6302);
      when "1100010011111" => q_unbuf <= my_rom(6303);
      when "1100010100000" => q_unbuf <= my_rom(6304);
      when "1100010100001" => q_unbuf <= my_rom(6305);
      when "1100010100010" => q_unbuf <= my_rom(6306);
      when "1100010100011" => q_unbuf <= my_rom(6307);
      when "1100010100100" => q_unbuf <= my_rom(6308);
      when "1100010100101" => q_unbuf <= my_rom(6309);
      when "1100010100110" => q_unbuf <= my_rom(6310);
      when "1100010100111" => q_unbuf <= my_rom(6311);
      when "1100010101000" => q_unbuf <= my_rom(6312);
      when "1100010101001" => q_unbuf <= my_rom(6313);
      when "1100010101010" => q_unbuf <= my_rom(6314);
      when "1100010101011" => q_unbuf <= my_rom(6315);
      when "1100010101100" => q_unbuf <= my_rom(6316);
      when "1100010101101" => q_unbuf <= my_rom(6317);
      when "1100010101110" => q_unbuf <= my_rom(6318);
      when "1100010101111" => q_unbuf <= my_rom(6319);
      when "1100010110000" => q_unbuf <= my_rom(6320);
      when "1100010110001" => q_unbuf <= my_rom(6321);
      when "1100010110010" => q_unbuf <= my_rom(6322);
      when "1100010110011" => q_unbuf <= my_rom(6323);
      when "1100010110100" => q_unbuf <= my_rom(6324);
      when "1100010110101" => q_unbuf <= my_rom(6325);
      when "1100010110110" => q_unbuf <= my_rom(6326);
      when "1100010110111" => q_unbuf <= my_rom(6327);
      when "1100010111000" => q_unbuf <= my_rom(6328);
      when "1100010111001" => q_unbuf <= my_rom(6329);
      when "1100010111010" => q_unbuf <= my_rom(6330);
      when "1100010111011" => q_unbuf <= my_rom(6331);
      when "1100010111100" => q_unbuf <= my_rom(6332);
      when "1100010111101" => q_unbuf <= my_rom(6333);
      when "1100010111110" => q_unbuf <= my_rom(6334);
      when "1100010111111" => q_unbuf <= my_rom(6335);
      when "1100011000000" => q_unbuf <= my_rom(6336);
      when "1100011000001" => q_unbuf <= my_rom(6337);
      when "1100011000010" => q_unbuf <= my_rom(6338);
      when "1100011000011" => q_unbuf <= my_rom(6339);
      when "1100011000100" => q_unbuf <= my_rom(6340);
      when "1100011000101" => q_unbuf <= my_rom(6341);
      when "1100011000110" => q_unbuf <= my_rom(6342);
      when "1100011000111" => q_unbuf <= my_rom(6343);
      when "1100011001000" => q_unbuf <= my_rom(6344);
      when "1100011001001" => q_unbuf <= my_rom(6345);
      when "1100011001010" => q_unbuf <= my_rom(6346);
      when "1100011001011" => q_unbuf <= my_rom(6347);
      when "1100011001100" => q_unbuf <= my_rom(6348);
      when "1100011001101" => q_unbuf <= my_rom(6349);
      when "1100011001110" => q_unbuf <= my_rom(6350);
      when "1100011001111" => q_unbuf <= my_rom(6351);
      when "1100011010000" => q_unbuf <= my_rom(6352);
      when "1100011010001" => q_unbuf <= my_rom(6353);
      when "1100011010010" => q_unbuf <= my_rom(6354);
      when "1100011010011" => q_unbuf <= my_rom(6355);
      when "1100011010100" => q_unbuf <= my_rom(6356);
      when "1100011010101" => q_unbuf <= my_rom(6357);
      when "1100011010110" => q_unbuf <= my_rom(6358);
      when "1100011010111" => q_unbuf <= my_rom(6359);
      when "1100011011000" => q_unbuf <= my_rom(6360);
      when "1100011011001" => q_unbuf <= my_rom(6361);
      when "1100011011010" => q_unbuf <= my_rom(6362);
      when "1100011011011" => q_unbuf <= my_rom(6363);
      when "1100011011100" => q_unbuf <= my_rom(6364);
      when "1100011011101" => q_unbuf <= my_rom(6365);
      when "1100011011110" => q_unbuf <= my_rom(6366);
      when "1100011011111" => q_unbuf <= my_rom(6367);
      when "1100011100000" => q_unbuf <= my_rom(6368);
      when "1100011100001" => q_unbuf <= my_rom(6369);
      when "1100011100010" => q_unbuf <= my_rom(6370);
      when "1100011100011" => q_unbuf <= my_rom(6371);
      when "1100011100100" => q_unbuf <= my_rom(6372);
      when "1100011100101" => q_unbuf <= my_rom(6373);
      when "1100011100110" => q_unbuf <= my_rom(6374);
      when "1100011100111" => q_unbuf <= my_rom(6375);
      when "1100011101000" => q_unbuf <= my_rom(6376);
      when "1100011101001" => q_unbuf <= my_rom(6377);
      when "1100011101010" => q_unbuf <= my_rom(6378);
      when "1100011101011" => q_unbuf <= my_rom(6379);
      when "1100011101100" => q_unbuf <= my_rom(6380);
      when "1100011101101" => q_unbuf <= my_rom(6381);
      when "1100011101110" => q_unbuf <= my_rom(6382);
      when "1100011101111" => q_unbuf <= my_rom(6383);
      when "1100011110000" => q_unbuf <= my_rom(6384);
      when "1100011110001" => q_unbuf <= my_rom(6385);
      when "1100011110010" => q_unbuf <= my_rom(6386);
      when "1100011110011" => q_unbuf <= my_rom(6387);
      when "1100011110100" => q_unbuf <= my_rom(6388);
      when "1100011110101" => q_unbuf <= my_rom(6389);
      when "1100011110110" => q_unbuf <= my_rom(6390);
      when "1100011110111" => q_unbuf <= my_rom(6391);
      when "1100011111000" => q_unbuf <= my_rom(6392);
      when "1100011111001" => q_unbuf <= my_rom(6393);
      when "1100011111010" => q_unbuf <= my_rom(6394);
      when "1100011111011" => q_unbuf <= my_rom(6395);
      when "1100011111100" => q_unbuf <= my_rom(6396);
      when "1100011111101" => q_unbuf <= my_rom(6397);
      when "1100011111110" => q_unbuf <= my_rom(6398);
      when "1100011111111" => q_unbuf <= my_rom(6399);
      when "1100100000000" => q_unbuf <= my_rom(6400);
      when "1100100000001" => q_unbuf <= my_rom(6401);
      when "1100100000010" => q_unbuf <= my_rom(6402);
      when "1100100000011" => q_unbuf <= my_rom(6403);
      when "1100100000100" => q_unbuf <= my_rom(6404);
      when "1100100000101" => q_unbuf <= my_rom(6405);
      when "1100100000110" => q_unbuf <= my_rom(6406);
      when "1100100000111" => q_unbuf <= my_rom(6407);
      when "1100100001000" => q_unbuf <= my_rom(6408);
      when "1100100001001" => q_unbuf <= my_rom(6409);
      when "1100100001010" => q_unbuf <= my_rom(6410);
      when "1100100001011" => q_unbuf <= my_rom(6411);
      when "1100100001100" => q_unbuf <= my_rom(6412);
      when "1100100001101" => q_unbuf <= my_rom(6413);
      when "1100100001110" => q_unbuf <= my_rom(6414);
      when "1100100001111" => q_unbuf <= my_rom(6415);
      when "1100100010000" => q_unbuf <= my_rom(6416);
      when "1100100010001" => q_unbuf <= my_rom(6417);
      when "1100100010010" => q_unbuf <= my_rom(6418);
      when "1100100010011" => q_unbuf <= my_rom(6419);
      when "1100100010100" => q_unbuf <= my_rom(6420);
      when "1100100010101" => q_unbuf <= my_rom(6421);
      when "1100100010110" => q_unbuf <= my_rom(6422);
      when "1100100010111" => q_unbuf <= my_rom(6423);
      when "1100100011000" => q_unbuf <= my_rom(6424);
      when "1100100011001" => q_unbuf <= my_rom(6425);
      when "1100100011010" => q_unbuf <= my_rom(6426);
      when "1100100011011" => q_unbuf <= my_rom(6427);
      when "1100100011100" => q_unbuf <= my_rom(6428);
      when "1100100011101" => q_unbuf <= my_rom(6429);
      when "1100100011110" => q_unbuf <= my_rom(6430);
      when "1100100011111" => q_unbuf <= my_rom(6431);
      when "1100100100000" => q_unbuf <= my_rom(6432);
      when "1100100100001" => q_unbuf <= my_rom(6433);
      when "1100100100010" => q_unbuf <= my_rom(6434);
      when "1100100100011" => q_unbuf <= my_rom(6435);
      when "1100100100100" => q_unbuf <= my_rom(6436);
      when "1100100100101" => q_unbuf <= my_rom(6437);
      when "1100100100110" => q_unbuf <= my_rom(6438);
      when "1100100100111" => q_unbuf <= my_rom(6439);
      when "1100100101000" => q_unbuf <= my_rom(6440);
      when "1100100101001" => q_unbuf <= my_rom(6441);
      when "1100100101010" => q_unbuf <= my_rom(6442);
      when "1100100101011" => q_unbuf <= my_rom(6443);
      when "1100100101100" => q_unbuf <= my_rom(6444);
      when "1100100101101" => q_unbuf <= my_rom(6445);
      when "1100100101110" => q_unbuf <= my_rom(6446);
      when "1100100101111" => q_unbuf <= my_rom(6447);
      when "1100100110000" => q_unbuf <= my_rom(6448);
      when "1100100110001" => q_unbuf <= my_rom(6449);
      when "1100100110010" => q_unbuf <= my_rom(6450);
      when "1100100110011" => q_unbuf <= my_rom(6451);
      when "1100100110100" => q_unbuf <= my_rom(6452);
      when "1100100110101" => q_unbuf <= my_rom(6453);
      when "1100100110110" => q_unbuf <= my_rom(6454);
      when "1100100110111" => q_unbuf <= my_rom(6455);
      when "1100100111000" => q_unbuf <= my_rom(6456);
      when "1100100111001" => q_unbuf <= my_rom(6457);
      when "1100100111010" => q_unbuf <= my_rom(6458);
      when "1100100111011" => q_unbuf <= my_rom(6459);
      when "1100100111100" => q_unbuf <= my_rom(6460);
      when "1100100111101" => q_unbuf <= my_rom(6461);
      when "1100100111110" => q_unbuf <= my_rom(6462);
      when "1100100111111" => q_unbuf <= my_rom(6463);
      when "1100101000000" => q_unbuf <= my_rom(6464);
      when "1100101000001" => q_unbuf <= my_rom(6465);
      when "1100101000010" => q_unbuf <= my_rom(6466);
      when "1100101000011" => q_unbuf <= my_rom(6467);
      when "1100101000100" => q_unbuf <= my_rom(6468);
      when "1100101000101" => q_unbuf <= my_rom(6469);
      when "1100101000110" => q_unbuf <= my_rom(6470);
      when "1100101000111" => q_unbuf <= my_rom(6471);
      when "1100101001000" => q_unbuf <= my_rom(6472);
      when "1100101001001" => q_unbuf <= my_rom(6473);
      when "1100101001010" => q_unbuf <= my_rom(6474);
      when "1100101001011" => q_unbuf <= my_rom(6475);
      when "1100101001100" => q_unbuf <= my_rom(6476);
      when "1100101001101" => q_unbuf <= my_rom(6477);
      when "1100101001110" => q_unbuf <= my_rom(6478);
      when "1100101001111" => q_unbuf <= my_rom(6479);
      when "1100101010000" => q_unbuf <= my_rom(6480);
      when "1100101010001" => q_unbuf <= my_rom(6481);
      when "1100101010010" => q_unbuf <= my_rom(6482);
      when "1100101010011" => q_unbuf <= my_rom(6483);
      when "1100101010100" => q_unbuf <= my_rom(6484);
      when "1100101010101" => q_unbuf <= my_rom(6485);
      when "1100101010110" => q_unbuf <= my_rom(6486);
      when "1100101010111" => q_unbuf <= my_rom(6487);
      when "1100101011000" => q_unbuf <= my_rom(6488);
      when "1100101011001" => q_unbuf <= my_rom(6489);
      when "1100101011010" => q_unbuf <= my_rom(6490);
      when "1100101011011" => q_unbuf <= my_rom(6491);
      when "1100101011100" => q_unbuf <= my_rom(6492);
      when "1100101011101" => q_unbuf <= my_rom(6493);
      when "1100101011110" => q_unbuf <= my_rom(6494);
      when "1100101011111" => q_unbuf <= my_rom(6495);
      when "1100101100000" => q_unbuf <= my_rom(6496);
      when "1100101100001" => q_unbuf <= my_rom(6497);
      when "1100101100010" => q_unbuf <= my_rom(6498);
      when "1100101100011" => q_unbuf <= my_rom(6499);
      when "1100101100100" => q_unbuf <= my_rom(6500);
      when "1100101100101" => q_unbuf <= my_rom(6501);
      when "1100101100110" => q_unbuf <= my_rom(6502);
      when "1100101100111" => q_unbuf <= my_rom(6503);
      when "1100101101000" => q_unbuf <= my_rom(6504);
      when "1100101101001" => q_unbuf <= my_rom(6505);
      when "1100101101010" => q_unbuf <= my_rom(6506);
      when "1100101101011" => q_unbuf <= my_rom(6507);
      when "1100101101100" => q_unbuf <= my_rom(6508);
      when "1100101101101" => q_unbuf <= my_rom(6509);
      when "1100101101110" => q_unbuf <= my_rom(6510);
      when "1100101101111" => q_unbuf <= my_rom(6511);
      when "1100101110000" => q_unbuf <= my_rom(6512);
      when "1100101110001" => q_unbuf <= my_rom(6513);
      when "1100101110010" => q_unbuf <= my_rom(6514);
      when "1100101110011" => q_unbuf <= my_rom(6515);
      when "1100101110100" => q_unbuf <= my_rom(6516);
      when "1100101110101" => q_unbuf <= my_rom(6517);
      when "1100101110110" => q_unbuf <= my_rom(6518);
      when "1100101110111" => q_unbuf <= my_rom(6519);
      when "1100101111000" => q_unbuf <= my_rom(6520);
      when "1100101111001" => q_unbuf <= my_rom(6521);
      when "1100101111010" => q_unbuf <= my_rom(6522);
      when "1100101111011" => q_unbuf <= my_rom(6523);
      when "1100101111100" => q_unbuf <= my_rom(6524);
      when "1100101111101" => q_unbuf <= my_rom(6525);
      when "1100101111110" => q_unbuf <= my_rom(6526);
      when "1100101111111" => q_unbuf <= my_rom(6527);
      when "1100110000000" => q_unbuf <= my_rom(6528);
      when "1100110000001" => q_unbuf <= my_rom(6529);
      when "1100110000010" => q_unbuf <= my_rom(6530);
      when "1100110000011" => q_unbuf <= my_rom(6531);
      when "1100110000100" => q_unbuf <= my_rom(6532);
      when "1100110000101" => q_unbuf <= my_rom(6533);
      when "1100110000110" => q_unbuf <= my_rom(6534);
      when "1100110000111" => q_unbuf <= my_rom(6535);
      when "1100110001000" => q_unbuf <= my_rom(6536);
      when "1100110001001" => q_unbuf <= my_rom(6537);
      when "1100110001010" => q_unbuf <= my_rom(6538);
      when "1100110001011" => q_unbuf <= my_rom(6539);
      when "1100110001100" => q_unbuf <= my_rom(6540);
      when "1100110001101" => q_unbuf <= my_rom(6541);
      when "1100110001110" => q_unbuf <= my_rom(6542);
      when "1100110001111" => q_unbuf <= my_rom(6543);
      when "1100110010000" => q_unbuf <= my_rom(6544);
      when "1100110010001" => q_unbuf <= my_rom(6545);
      when "1100110010010" => q_unbuf <= my_rom(6546);
      when "1100110010011" => q_unbuf <= my_rom(6547);
      when "1100110010100" => q_unbuf <= my_rom(6548);
      when "1100110010101" => q_unbuf <= my_rom(6549);
      when "1100110010110" => q_unbuf <= my_rom(6550);
      when "1100110010111" => q_unbuf <= my_rom(6551);
      when "1100110011000" => q_unbuf <= my_rom(6552);
      when "1100110011001" => q_unbuf <= my_rom(6553);
      when "1100110011010" => q_unbuf <= my_rom(6554);
      when "1100110011011" => q_unbuf <= my_rom(6555);
      when "1100110011100" => q_unbuf <= my_rom(6556);
      when "1100110011101" => q_unbuf <= my_rom(6557);
      when "1100110011110" => q_unbuf <= my_rom(6558);
      when "1100110011111" => q_unbuf <= my_rom(6559);
      when "1100110100000" => q_unbuf <= my_rom(6560);
      when "1100110100001" => q_unbuf <= my_rom(6561);
      when "1100110100010" => q_unbuf <= my_rom(6562);
      when "1100110100011" => q_unbuf <= my_rom(6563);
      when "1100110100100" => q_unbuf <= my_rom(6564);
      when "1100110100101" => q_unbuf <= my_rom(6565);
      when "1100110100110" => q_unbuf <= my_rom(6566);
      when "1100110100111" => q_unbuf <= my_rom(6567);
      when "1100110101000" => q_unbuf <= my_rom(6568);
      when "1100110101001" => q_unbuf <= my_rom(6569);
      when "1100110101010" => q_unbuf <= my_rom(6570);
      when "1100110101011" => q_unbuf <= my_rom(6571);
      when "1100110101100" => q_unbuf <= my_rom(6572);
      when "1100110101101" => q_unbuf <= my_rom(6573);
      when "1100110101110" => q_unbuf <= my_rom(6574);
      when "1100110101111" => q_unbuf <= my_rom(6575);
      when "1100110110000" => q_unbuf <= my_rom(6576);
      when "1100110110001" => q_unbuf <= my_rom(6577);
      when "1100110110010" => q_unbuf <= my_rom(6578);
      when "1100110110011" => q_unbuf <= my_rom(6579);
      when "1100110110100" => q_unbuf <= my_rom(6580);
      when "1100110110101" => q_unbuf <= my_rom(6581);
      when "1100110110110" => q_unbuf <= my_rom(6582);
      when "1100110110111" => q_unbuf <= my_rom(6583);
      when "1100110111000" => q_unbuf <= my_rom(6584);
      when "1100110111001" => q_unbuf <= my_rom(6585);
      when "1100110111010" => q_unbuf <= my_rom(6586);
      when "1100110111011" => q_unbuf <= my_rom(6587);
      when "1100110111100" => q_unbuf <= my_rom(6588);
      when "1100110111101" => q_unbuf <= my_rom(6589);
      when "1100110111110" => q_unbuf <= my_rom(6590);
      when "1100110111111" => q_unbuf <= my_rom(6591);
      when "1100111000000" => q_unbuf <= my_rom(6592);
      when "1100111000001" => q_unbuf <= my_rom(6593);
      when "1100111000010" => q_unbuf <= my_rom(6594);
      when "1100111000011" => q_unbuf <= my_rom(6595);
      when "1100111000100" => q_unbuf <= my_rom(6596);
      when "1100111000101" => q_unbuf <= my_rom(6597);
      when "1100111000110" => q_unbuf <= my_rom(6598);
      when "1100111000111" => q_unbuf <= my_rom(6599);
      when "1100111001000" => q_unbuf <= my_rom(6600);
      when "1100111001001" => q_unbuf <= my_rom(6601);
      when "1100111001010" => q_unbuf <= my_rom(6602);
      when "1100111001011" => q_unbuf <= my_rom(6603);
      when "1100111001100" => q_unbuf <= my_rom(6604);
      when "1100111001101" => q_unbuf <= my_rom(6605);
      when "1100111001110" => q_unbuf <= my_rom(6606);
      when "1100111001111" => q_unbuf <= my_rom(6607);
      when "1100111010000" => q_unbuf <= my_rom(6608);
      when "1100111010001" => q_unbuf <= my_rom(6609);
      when "1100111010010" => q_unbuf <= my_rom(6610);
      when "1100111010011" => q_unbuf <= my_rom(6611);
      when "1100111010100" => q_unbuf <= my_rom(6612);
      when "1100111010101" => q_unbuf <= my_rom(6613);
      when "1100111010110" => q_unbuf <= my_rom(6614);
      when "1100111010111" => q_unbuf <= my_rom(6615);
      when "1100111011000" => q_unbuf <= my_rom(6616);
      when "1100111011001" => q_unbuf <= my_rom(6617);
      when "1100111011010" => q_unbuf <= my_rom(6618);
      when "1100111011011" => q_unbuf <= my_rom(6619);
      when "1100111011100" => q_unbuf <= my_rom(6620);
      when "1100111011101" => q_unbuf <= my_rom(6621);
      when "1100111011110" => q_unbuf <= my_rom(6622);
      when "1100111011111" => q_unbuf <= my_rom(6623);
      when "1100111100000" => q_unbuf <= my_rom(6624);
      when "1100111100001" => q_unbuf <= my_rom(6625);
      when "1100111100010" => q_unbuf <= my_rom(6626);
      when "1100111100011" => q_unbuf <= my_rom(6627);
      when "1100111100100" => q_unbuf <= my_rom(6628);
      when "1100111100101" => q_unbuf <= my_rom(6629);
      when "1100111100110" => q_unbuf <= my_rom(6630);
      when "1100111100111" => q_unbuf <= my_rom(6631);
      when "1100111101000" => q_unbuf <= my_rom(6632);
      when "1100111101001" => q_unbuf <= my_rom(6633);
      when "1100111101010" => q_unbuf <= my_rom(6634);
      when "1100111101011" => q_unbuf <= my_rom(6635);
      when "1100111101100" => q_unbuf <= my_rom(6636);
      when "1100111101101" => q_unbuf <= my_rom(6637);
      when "1100111101110" => q_unbuf <= my_rom(6638);
      when "1100111101111" => q_unbuf <= my_rom(6639);
      when "1100111110000" => q_unbuf <= my_rom(6640);
      when "1100111110001" => q_unbuf <= my_rom(6641);
      when "1100111110010" => q_unbuf <= my_rom(6642);
      when "1100111110011" => q_unbuf <= my_rom(6643);
      when "1100111110100" => q_unbuf <= my_rom(6644);
      when "1100111110101" => q_unbuf <= my_rom(6645);
      when "1100111110110" => q_unbuf <= my_rom(6646);
      when "1100111110111" => q_unbuf <= my_rom(6647);
      when "1100111111000" => q_unbuf <= my_rom(6648);
      when "1100111111001" => q_unbuf <= my_rom(6649);
      when "1100111111010" => q_unbuf <= my_rom(6650);
      when "1100111111011" => q_unbuf <= my_rom(6651);
      when "1100111111100" => q_unbuf <= my_rom(6652);
      when "1100111111101" => q_unbuf <= my_rom(6653);
      when "1100111111110" => q_unbuf <= my_rom(6654);
      when "1100111111111" => q_unbuf <= my_rom(6655);
      when "1101000000000" => q_unbuf <= my_rom(6656);
      when "1101000000001" => q_unbuf <= my_rom(6657);
      when "1101000000010" => q_unbuf <= my_rom(6658);
      when "1101000000011" => q_unbuf <= my_rom(6659);
      when "1101000000100" => q_unbuf <= my_rom(6660);
      when "1101000000101" => q_unbuf <= my_rom(6661);
      when "1101000000110" => q_unbuf <= my_rom(6662);
      when "1101000000111" => q_unbuf <= my_rom(6663);
      when "1101000001000" => q_unbuf <= my_rom(6664);
      when "1101000001001" => q_unbuf <= my_rom(6665);
      when "1101000001010" => q_unbuf <= my_rom(6666);
      when "1101000001011" => q_unbuf <= my_rom(6667);
      when "1101000001100" => q_unbuf <= my_rom(6668);
      when "1101000001101" => q_unbuf <= my_rom(6669);
      when "1101000001110" => q_unbuf <= my_rom(6670);
      when "1101000001111" => q_unbuf <= my_rom(6671);
      when "1101000010000" => q_unbuf <= my_rom(6672);
      when "1101000010001" => q_unbuf <= my_rom(6673);
      when "1101000010010" => q_unbuf <= my_rom(6674);
      when "1101000010011" => q_unbuf <= my_rom(6675);
      when "1101000010100" => q_unbuf <= my_rom(6676);
      when "1101000010101" => q_unbuf <= my_rom(6677);
      when "1101000010110" => q_unbuf <= my_rom(6678);
      when "1101000010111" => q_unbuf <= my_rom(6679);
      when "1101000011000" => q_unbuf <= my_rom(6680);
      when "1101000011001" => q_unbuf <= my_rom(6681);
      when "1101000011010" => q_unbuf <= my_rom(6682);
      when "1101000011011" => q_unbuf <= my_rom(6683);
      when "1101000011100" => q_unbuf <= my_rom(6684);
      when "1101000011101" => q_unbuf <= my_rom(6685);
      when "1101000011110" => q_unbuf <= my_rom(6686);
      when "1101000011111" => q_unbuf <= my_rom(6687);
      when "1101000100000" => q_unbuf <= my_rom(6688);
      when "1101000100001" => q_unbuf <= my_rom(6689);
      when "1101000100010" => q_unbuf <= my_rom(6690);
      when "1101000100011" => q_unbuf <= my_rom(6691);
      when "1101000100100" => q_unbuf <= my_rom(6692);
      when "1101000100101" => q_unbuf <= my_rom(6693);
      when "1101000100110" => q_unbuf <= my_rom(6694);
      when "1101000100111" => q_unbuf <= my_rom(6695);
      when "1101000101000" => q_unbuf <= my_rom(6696);
      when "1101000101001" => q_unbuf <= my_rom(6697);
      when "1101000101010" => q_unbuf <= my_rom(6698);
      when "1101000101011" => q_unbuf <= my_rom(6699);
      when "1101000101100" => q_unbuf <= my_rom(6700);
      when "1101000101101" => q_unbuf <= my_rom(6701);
      when "1101000101110" => q_unbuf <= my_rom(6702);
      when "1101000101111" => q_unbuf <= my_rom(6703);
      when "1101000110000" => q_unbuf <= my_rom(6704);
      when "1101000110001" => q_unbuf <= my_rom(6705);
      when "1101000110010" => q_unbuf <= my_rom(6706);
      when "1101000110011" => q_unbuf <= my_rom(6707);
      when "1101000110100" => q_unbuf <= my_rom(6708);
      when "1101000110101" => q_unbuf <= my_rom(6709);
      when "1101000110110" => q_unbuf <= my_rom(6710);
      when "1101000110111" => q_unbuf <= my_rom(6711);
      when "1101000111000" => q_unbuf <= my_rom(6712);
      when "1101000111001" => q_unbuf <= my_rom(6713);
      when "1101000111010" => q_unbuf <= my_rom(6714);
      when "1101000111011" => q_unbuf <= my_rom(6715);
      when "1101000111100" => q_unbuf <= my_rom(6716);
      when "1101000111101" => q_unbuf <= my_rom(6717);
      when "1101000111110" => q_unbuf <= my_rom(6718);
      when "1101000111111" => q_unbuf <= my_rom(6719);
      when "1101001000000" => q_unbuf <= my_rom(6720);
      when "1101001000001" => q_unbuf <= my_rom(6721);
      when "1101001000010" => q_unbuf <= my_rom(6722);
      when "1101001000011" => q_unbuf <= my_rom(6723);
      when "1101001000100" => q_unbuf <= my_rom(6724);
      when "1101001000101" => q_unbuf <= my_rom(6725);
      when "1101001000110" => q_unbuf <= my_rom(6726);
      when "1101001000111" => q_unbuf <= my_rom(6727);
      when "1101001001000" => q_unbuf <= my_rom(6728);
      when "1101001001001" => q_unbuf <= my_rom(6729);
      when "1101001001010" => q_unbuf <= my_rom(6730);
      when "1101001001011" => q_unbuf <= my_rom(6731);
      when "1101001001100" => q_unbuf <= my_rom(6732);
      when "1101001001101" => q_unbuf <= my_rom(6733);
      when "1101001001110" => q_unbuf <= my_rom(6734);
      when "1101001001111" => q_unbuf <= my_rom(6735);
      when "1101001010000" => q_unbuf <= my_rom(6736);
      when "1101001010001" => q_unbuf <= my_rom(6737);
      when "1101001010010" => q_unbuf <= my_rom(6738);
      when "1101001010011" => q_unbuf <= my_rom(6739);
      when "1101001010100" => q_unbuf <= my_rom(6740);
      when "1101001010101" => q_unbuf <= my_rom(6741);
      when "1101001010110" => q_unbuf <= my_rom(6742);
      when "1101001010111" => q_unbuf <= my_rom(6743);
      when "1101001011000" => q_unbuf <= my_rom(6744);
      when "1101001011001" => q_unbuf <= my_rom(6745);
      when "1101001011010" => q_unbuf <= my_rom(6746);
      when "1101001011011" => q_unbuf <= my_rom(6747);
      when "1101001011100" => q_unbuf <= my_rom(6748);
      when "1101001011101" => q_unbuf <= my_rom(6749);
      when "1101001011110" => q_unbuf <= my_rom(6750);
      when "1101001011111" => q_unbuf <= my_rom(6751);
      when "1101001100000" => q_unbuf <= my_rom(6752);
      when "1101001100001" => q_unbuf <= my_rom(6753);
      when "1101001100010" => q_unbuf <= my_rom(6754);
      when "1101001100011" => q_unbuf <= my_rom(6755);
      when "1101001100100" => q_unbuf <= my_rom(6756);
      when "1101001100101" => q_unbuf <= my_rom(6757);
      when "1101001100110" => q_unbuf <= my_rom(6758);
      when "1101001100111" => q_unbuf <= my_rom(6759);
      when "1101001101000" => q_unbuf <= my_rom(6760);
      when "1101001101001" => q_unbuf <= my_rom(6761);
      when "1101001101010" => q_unbuf <= my_rom(6762);
      when "1101001101011" => q_unbuf <= my_rom(6763);
      when "1101001101100" => q_unbuf <= my_rom(6764);
      when "1101001101101" => q_unbuf <= my_rom(6765);
      when "1101001101110" => q_unbuf <= my_rom(6766);
      when "1101001101111" => q_unbuf <= my_rom(6767);
      when "1101001110000" => q_unbuf <= my_rom(6768);
      when "1101001110001" => q_unbuf <= my_rom(6769);
      when "1101001110010" => q_unbuf <= my_rom(6770);
      when "1101001110011" => q_unbuf <= my_rom(6771);
      when "1101001110100" => q_unbuf <= my_rom(6772);
      when "1101001110101" => q_unbuf <= my_rom(6773);
      when "1101001110110" => q_unbuf <= my_rom(6774);
      when "1101001110111" => q_unbuf <= my_rom(6775);
      when "1101001111000" => q_unbuf <= my_rom(6776);
      when "1101001111001" => q_unbuf <= my_rom(6777);
      when "1101001111010" => q_unbuf <= my_rom(6778);
      when "1101001111011" => q_unbuf <= my_rom(6779);
      when "1101001111100" => q_unbuf <= my_rom(6780);
      when "1101001111101" => q_unbuf <= my_rom(6781);
      when "1101001111110" => q_unbuf <= my_rom(6782);
      when "1101001111111" => q_unbuf <= my_rom(6783);
      when "1101010000000" => q_unbuf <= my_rom(6784);
      when "1101010000001" => q_unbuf <= my_rom(6785);
      when "1101010000010" => q_unbuf <= my_rom(6786);
      when "1101010000011" => q_unbuf <= my_rom(6787);
      when "1101010000100" => q_unbuf <= my_rom(6788);
      when "1101010000101" => q_unbuf <= my_rom(6789);
      when "1101010000110" => q_unbuf <= my_rom(6790);
      when "1101010000111" => q_unbuf <= my_rom(6791);
      when "1101010001000" => q_unbuf <= my_rom(6792);
      when "1101010001001" => q_unbuf <= my_rom(6793);
      when "1101010001010" => q_unbuf <= my_rom(6794);
      when "1101010001011" => q_unbuf <= my_rom(6795);
      when "1101010001100" => q_unbuf <= my_rom(6796);
      when "1101010001101" => q_unbuf <= my_rom(6797);
      when "1101010001110" => q_unbuf <= my_rom(6798);
      when "1101010001111" => q_unbuf <= my_rom(6799);
      when "1101010010000" => q_unbuf <= my_rom(6800);
      when "1101010010001" => q_unbuf <= my_rom(6801);
      when "1101010010010" => q_unbuf <= my_rom(6802);
      when "1101010010011" => q_unbuf <= my_rom(6803);
      when "1101010010100" => q_unbuf <= my_rom(6804);
      when "1101010010101" => q_unbuf <= my_rom(6805);
      when "1101010010110" => q_unbuf <= my_rom(6806);
      when "1101010010111" => q_unbuf <= my_rom(6807);
      when "1101010011000" => q_unbuf <= my_rom(6808);
      when "1101010011001" => q_unbuf <= my_rom(6809);
      when "1101010011010" => q_unbuf <= my_rom(6810);
      when "1101010011011" => q_unbuf <= my_rom(6811);
      when "1101010011100" => q_unbuf <= my_rom(6812);
      when "1101010011101" => q_unbuf <= my_rom(6813);
      when "1101010011110" => q_unbuf <= my_rom(6814);
      when "1101010011111" => q_unbuf <= my_rom(6815);
      when "1101010100000" => q_unbuf <= my_rom(6816);
      when "1101010100001" => q_unbuf <= my_rom(6817);
      when "1101010100010" => q_unbuf <= my_rom(6818);
      when "1101010100011" => q_unbuf <= my_rom(6819);
      when "1101010100100" => q_unbuf <= my_rom(6820);
      when "1101010100101" => q_unbuf <= my_rom(6821);
      when "1101010100110" => q_unbuf <= my_rom(6822);
      when "1101010100111" => q_unbuf <= my_rom(6823);
      when "1101010101000" => q_unbuf <= my_rom(6824);
      when "1101010101001" => q_unbuf <= my_rom(6825);
      when "1101010101010" => q_unbuf <= my_rom(6826);
      when "1101010101011" => q_unbuf <= my_rom(6827);
      when "1101010101100" => q_unbuf <= my_rom(6828);
      when "1101010101101" => q_unbuf <= my_rom(6829);
      when "1101010101110" => q_unbuf <= my_rom(6830);
      when "1101010101111" => q_unbuf <= my_rom(6831);
      when "1101010110000" => q_unbuf <= my_rom(6832);
      when "1101010110001" => q_unbuf <= my_rom(6833);
      when "1101010110010" => q_unbuf <= my_rom(6834);
      when "1101010110011" => q_unbuf <= my_rom(6835);
      when "1101010110100" => q_unbuf <= my_rom(6836);
      when "1101010110101" => q_unbuf <= my_rom(6837);
      when "1101010110110" => q_unbuf <= my_rom(6838);
      when "1101010110111" => q_unbuf <= my_rom(6839);
      when "1101010111000" => q_unbuf <= my_rom(6840);
      when "1101010111001" => q_unbuf <= my_rom(6841);
      when "1101010111010" => q_unbuf <= my_rom(6842);
      when "1101010111011" => q_unbuf <= my_rom(6843);
      when "1101010111100" => q_unbuf <= my_rom(6844);
      when "1101010111101" => q_unbuf <= my_rom(6845);
      when "1101010111110" => q_unbuf <= my_rom(6846);
      when "1101010111111" => q_unbuf <= my_rom(6847);
      when "1101011000000" => q_unbuf <= my_rom(6848);
      when "1101011000001" => q_unbuf <= my_rom(6849);
      when "1101011000010" => q_unbuf <= my_rom(6850);
      when "1101011000011" => q_unbuf <= my_rom(6851);
      when "1101011000100" => q_unbuf <= my_rom(6852);
      when "1101011000101" => q_unbuf <= my_rom(6853);
      when "1101011000110" => q_unbuf <= my_rom(6854);
      when "1101011000111" => q_unbuf <= my_rom(6855);
      when "1101011001000" => q_unbuf <= my_rom(6856);
      when "1101011001001" => q_unbuf <= my_rom(6857);
      when "1101011001010" => q_unbuf <= my_rom(6858);
      when "1101011001011" => q_unbuf <= my_rom(6859);
      when "1101011001100" => q_unbuf <= my_rom(6860);
      when "1101011001101" => q_unbuf <= my_rom(6861);
      when "1101011001110" => q_unbuf <= my_rom(6862);
      when "1101011001111" => q_unbuf <= my_rom(6863);
      when "1101011010000" => q_unbuf <= my_rom(6864);
      when "1101011010001" => q_unbuf <= my_rom(6865);
      when "1101011010010" => q_unbuf <= my_rom(6866);
      when "1101011010011" => q_unbuf <= my_rom(6867);
      when "1101011010100" => q_unbuf <= my_rom(6868);
      when "1101011010101" => q_unbuf <= my_rom(6869);
      when "1101011010110" => q_unbuf <= my_rom(6870);
      when "1101011010111" => q_unbuf <= my_rom(6871);
      when "1101011011000" => q_unbuf <= my_rom(6872);
      when "1101011011001" => q_unbuf <= my_rom(6873);
      when "1101011011010" => q_unbuf <= my_rom(6874);
      when "1101011011011" => q_unbuf <= my_rom(6875);
      when "1101011011100" => q_unbuf <= my_rom(6876);
      when "1101011011101" => q_unbuf <= my_rom(6877);
      when "1101011011110" => q_unbuf <= my_rom(6878);
      when "1101011011111" => q_unbuf <= my_rom(6879);
      when "1101011100000" => q_unbuf <= my_rom(6880);
      when "1101011100001" => q_unbuf <= my_rom(6881);
      when "1101011100010" => q_unbuf <= my_rom(6882);
      when "1101011100011" => q_unbuf <= my_rom(6883);
      when "1101011100100" => q_unbuf <= my_rom(6884);
      when "1101011100101" => q_unbuf <= my_rom(6885);
      when "1101011100110" => q_unbuf <= my_rom(6886);
      when "1101011100111" => q_unbuf <= my_rom(6887);
      when "1101011101000" => q_unbuf <= my_rom(6888);
      when "1101011101001" => q_unbuf <= my_rom(6889);
      when "1101011101010" => q_unbuf <= my_rom(6890);
      when "1101011101011" => q_unbuf <= my_rom(6891);
      when "1101011101100" => q_unbuf <= my_rom(6892);
      when "1101011101101" => q_unbuf <= my_rom(6893);
      when "1101011101110" => q_unbuf <= my_rom(6894);
      when "1101011101111" => q_unbuf <= my_rom(6895);
      when "1101011110000" => q_unbuf <= my_rom(6896);
      when "1101011110001" => q_unbuf <= my_rom(6897);
      when "1101011110010" => q_unbuf <= my_rom(6898);
      when "1101011110011" => q_unbuf <= my_rom(6899);
      when "1101011110100" => q_unbuf <= my_rom(6900);
      when "1101011110101" => q_unbuf <= my_rom(6901);
      when "1101011110110" => q_unbuf <= my_rom(6902);
      when "1101011110111" => q_unbuf <= my_rom(6903);
      when "1101011111000" => q_unbuf <= my_rom(6904);
      when "1101011111001" => q_unbuf <= my_rom(6905);
      when "1101011111010" => q_unbuf <= my_rom(6906);
      when "1101011111011" => q_unbuf <= my_rom(6907);
      when "1101011111100" => q_unbuf <= my_rom(6908);
      when "1101011111101" => q_unbuf <= my_rom(6909);
      when "1101011111110" => q_unbuf <= my_rom(6910);
      when "1101011111111" => q_unbuf <= my_rom(6911);
      when "1101100000000" => q_unbuf <= my_rom(6912);
      when "1101100000001" => q_unbuf <= my_rom(6913);
      when "1101100000010" => q_unbuf <= my_rom(6914);
      when "1101100000011" => q_unbuf <= my_rom(6915);
      when "1101100000100" => q_unbuf <= my_rom(6916);
      when "1101100000101" => q_unbuf <= my_rom(6917);
      when "1101100000110" => q_unbuf <= my_rom(6918);
      when "1101100000111" => q_unbuf <= my_rom(6919);
      when "1101100001000" => q_unbuf <= my_rom(6920);
      when "1101100001001" => q_unbuf <= my_rom(6921);
      when "1101100001010" => q_unbuf <= my_rom(6922);
      when "1101100001011" => q_unbuf <= my_rom(6923);
      when "1101100001100" => q_unbuf <= my_rom(6924);
      when "1101100001101" => q_unbuf <= my_rom(6925);
      when "1101100001110" => q_unbuf <= my_rom(6926);
      when "1101100001111" => q_unbuf <= my_rom(6927);
      when "1101100010000" => q_unbuf <= my_rom(6928);
      when "1101100010001" => q_unbuf <= my_rom(6929);
      when "1101100010010" => q_unbuf <= my_rom(6930);
      when "1101100010011" => q_unbuf <= my_rom(6931);
      when "1101100010100" => q_unbuf <= my_rom(6932);
      when "1101100010101" => q_unbuf <= my_rom(6933);
      when "1101100010110" => q_unbuf <= my_rom(6934);
      when "1101100010111" => q_unbuf <= my_rom(6935);
      when "1101100011000" => q_unbuf <= my_rom(6936);
      when "1101100011001" => q_unbuf <= my_rom(6937);
      when "1101100011010" => q_unbuf <= my_rom(6938);
      when "1101100011011" => q_unbuf <= my_rom(6939);
      when "1101100011100" => q_unbuf <= my_rom(6940);
      when "1101100011101" => q_unbuf <= my_rom(6941);
      when "1101100011110" => q_unbuf <= my_rom(6942);
      when "1101100011111" => q_unbuf <= my_rom(6943);
      when "1101100100000" => q_unbuf <= my_rom(6944);
      when "1101100100001" => q_unbuf <= my_rom(6945);
      when "1101100100010" => q_unbuf <= my_rom(6946);
      when "1101100100011" => q_unbuf <= my_rom(6947);
      when "1101100100100" => q_unbuf <= my_rom(6948);
      when "1101100100101" => q_unbuf <= my_rom(6949);
      when "1101100100110" => q_unbuf <= my_rom(6950);
      when "1101100100111" => q_unbuf <= my_rom(6951);
      when "1101100101000" => q_unbuf <= my_rom(6952);
      when "1101100101001" => q_unbuf <= my_rom(6953);
      when "1101100101010" => q_unbuf <= my_rom(6954);
      when "1101100101011" => q_unbuf <= my_rom(6955);
      when "1101100101100" => q_unbuf <= my_rom(6956);
      when "1101100101101" => q_unbuf <= my_rom(6957);
      when "1101100101110" => q_unbuf <= my_rom(6958);
      when "1101100101111" => q_unbuf <= my_rom(6959);
      when "1101100110000" => q_unbuf <= my_rom(6960);
      when "1101100110001" => q_unbuf <= my_rom(6961);
      when "1101100110010" => q_unbuf <= my_rom(6962);
      when "1101100110011" => q_unbuf <= my_rom(6963);
      when "1101100110100" => q_unbuf <= my_rom(6964);
      when "1101100110101" => q_unbuf <= my_rom(6965);
      when "1101100110110" => q_unbuf <= my_rom(6966);
      when "1101100110111" => q_unbuf <= my_rom(6967);
      when "1101100111000" => q_unbuf <= my_rom(6968);
      when "1101100111001" => q_unbuf <= my_rom(6969);
      when "1101100111010" => q_unbuf <= my_rom(6970);
      when "1101100111011" => q_unbuf <= my_rom(6971);
      when "1101100111100" => q_unbuf <= my_rom(6972);
      when "1101100111101" => q_unbuf <= my_rom(6973);
      when "1101100111110" => q_unbuf <= my_rom(6974);
      when "1101100111111" => q_unbuf <= my_rom(6975);
      when "1101101000000" => q_unbuf <= my_rom(6976);
      when "1101101000001" => q_unbuf <= my_rom(6977);
      when "1101101000010" => q_unbuf <= my_rom(6978);
      when "1101101000011" => q_unbuf <= my_rom(6979);
      when "1101101000100" => q_unbuf <= my_rom(6980);
      when "1101101000101" => q_unbuf <= my_rom(6981);
      when "1101101000110" => q_unbuf <= my_rom(6982);
      when "1101101000111" => q_unbuf <= my_rom(6983);
      when "1101101001000" => q_unbuf <= my_rom(6984);
      when "1101101001001" => q_unbuf <= my_rom(6985);
      when "1101101001010" => q_unbuf <= my_rom(6986);
      when "1101101001011" => q_unbuf <= my_rom(6987);
      when "1101101001100" => q_unbuf <= my_rom(6988);
      when "1101101001101" => q_unbuf <= my_rom(6989);
      when "1101101001110" => q_unbuf <= my_rom(6990);
      when "1101101001111" => q_unbuf <= my_rom(6991);
      when "1101101010000" => q_unbuf <= my_rom(6992);
      when "1101101010001" => q_unbuf <= my_rom(6993);
      when "1101101010010" => q_unbuf <= my_rom(6994);
      when "1101101010011" => q_unbuf <= my_rom(6995);
      when "1101101010100" => q_unbuf <= my_rom(6996);
      when "1101101010101" => q_unbuf <= my_rom(6997);
      when "1101101010110" => q_unbuf <= my_rom(6998);
      when "1101101010111" => q_unbuf <= my_rom(6999);
      when "1101101011000" => q_unbuf <= my_rom(7000);
      when "1101101011001" => q_unbuf <= my_rom(7001);
      when "1101101011010" => q_unbuf <= my_rom(7002);
      when "1101101011011" => q_unbuf <= my_rom(7003);
      when "1101101011100" => q_unbuf <= my_rom(7004);
      when "1101101011101" => q_unbuf <= my_rom(7005);
      when "1101101011110" => q_unbuf <= my_rom(7006);
      when "1101101011111" => q_unbuf <= my_rom(7007);
      when "1101101100000" => q_unbuf <= my_rom(7008);
      when "1101101100001" => q_unbuf <= my_rom(7009);
      when "1101101100010" => q_unbuf <= my_rom(7010);
      when "1101101100011" => q_unbuf <= my_rom(7011);
      when "1101101100100" => q_unbuf <= my_rom(7012);
      when "1101101100101" => q_unbuf <= my_rom(7013);
      when "1101101100110" => q_unbuf <= my_rom(7014);
      when "1101101100111" => q_unbuf <= my_rom(7015);
      when "1101101101000" => q_unbuf <= my_rom(7016);
      when "1101101101001" => q_unbuf <= my_rom(7017);
      when "1101101101010" => q_unbuf <= my_rom(7018);
      when "1101101101011" => q_unbuf <= my_rom(7019);
      when "1101101101100" => q_unbuf <= my_rom(7020);
      when "1101101101101" => q_unbuf <= my_rom(7021);
      when "1101101101110" => q_unbuf <= my_rom(7022);
      when "1101101101111" => q_unbuf <= my_rom(7023);
      when "1101101110000" => q_unbuf <= my_rom(7024);
      when "1101101110001" => q_unbuf <= my_rom(7025);
      when "1101101110010" => q_unbuf <= my_rom(7026);
      when "1101101110011" => q_unbuf <= my_rom(7027);
      when "1101101110100" => q_unbuf <= my_rom(7028);
      when "1101101110101" => q_unbuf <= my_rom(7029);
      when "1101101110110" => q_unbuf <= my_rom(7030);
      when "1101101110111" => q_unbuf <= my_rom(7031);
      when "1101101111000" => q_unbuf <= my_rom(7032);
      when "1101101111001" => q_unbuf <= my_rom(7033);
      when "1101101111010" => q_unbuf <= my_rom(7034);
      when "1101101111011" => q_unbuf <= my_rom(7035);
      when "1101101111100" => q_unbuf <= my_rom(7036);
      when "1101101111101" => q_unbuf <= my_rom(7037);
      when "1101101111110" => q_unbuf <= my_rom(7038);
      when "1101101111111" => q_unbuf <= my_rom(7039);
      when "1101110000000" => q_unbuf <= my_rom(7040);
      when "1101110000001" => q_unbuf <= my_rom(7041);
      when "1101110000010" => q_unbuf <= my_rom(7042);
      when "1101110000011" => q_unbuf <= my_rom(7043);
      when "1101110000100" => q_unbuf <= my_rom(7044);
      when "1101110000101" => q_unbuf <= my_rom(7045);
      when "1101110000110" => q_unbuf <= my_rom(7046);
      when "1101110000111" => q_unbuf <= my_rom(7047);
      when "1101110001000" => q_unbuf <= my_rom(7048);
      when "1101110001001" => q_unbuf <= my_rom(7049);
      when "1101110001010" => q_unbuf <= my_rom(7050);
      when "1101110001011" => q_unbuf <= my_rom(7051);
      when "1101110001100" => q_unbuf <= my_rom(7052);
      when "1101110001101" => q_unbuf <= my_rom(7053);
      when "1101110001110" => q_unbuf <= my_rom(7054);
      when "1101110001111" => q_unbuf <= my_rom(7055);
      when "1101110010000" => q_unbuf <= my_rom(7056);
      when "1101110010001" => q_unbuf <= my_rom(7057);
      when "1101110010010" => q_unbuf <= my_rom(7058);
      when "1101110010011" => q_unbuf <= my_rom(7059);
      when "1101110010100" => q_unbuf <= my_rom(7060);
      when "1101110010101" => q_unbuf <= my_rom(7061);
      when "1101110010110" => q_unbuf <= my_rom(7062);
      when "1101110010111" => q_unbuf <= my_rom(7063);
      when "1101110011000" => q_unbuf <= my_rom(7064);
      when "1101110011001" => q_unbuf <= my_rom(7065);
      when "1101110011010" => q_unbuf <= my_rom(7066);
      when "1101110011011" => q_unbuf <= my_rom(7067);
      when "1101110011100" => q_unbuf <= my_rom(7068);
      when "1101110011101" => q_unbuf <= my_rom(7069);
      when "1101110011110" => q_unbuf <= my_rom(7070);
      when "1101110011111" => q_unbuf <= my_rom(7071);
      when "1101110100000" => q_unbuf <= my_rom(7072);
      when "1101110100001" => q_unbuf <= my_rom(7073);
      when "1101110100010" => q_unbuf <= my_rom(7074);
      when "1101110100011" => q_unbuf <= my_rom(7075);
      when "1101110100100" => q_unbuf <= my_rom(7076);
      when "1101110100101" => q_unbuf <= my_rom(7077);
      when "1101110100110" => q_unbuf <= my_rom(7078);
      when "1101110100111" => q_unbuf <= my_rom(7079);
      when "1101110101000" => q_unbuf <= my_rom(7080);
      when "1101110101001" => q_unbuf <= my_rom(7081);
      when "1101110101010" => q_unbuf <= my_rom(7082);
      when "1101110101011" => q_unbuf <= my_rom(7083);
      when "1101110101100" => q_unbuf <= my_rom(7084);
      when "1101110101101" => q_unbuf <= my_rom(7085);
      when "1101110101110" => q_unbuf <= my_rom(7086);
      when "1101110101111" => q_unbuf <= my_rom(7087);
      when "1101110110000" => q_unbuf <= my_rom(7088);
      when "1101110110001" => q_unbuf <= my_rom(7089);
      when "1101110110010" => q_unbuf <= my_rom(7090);
      when "1101110110011" => q_unbuf <= my_rom(7091);
      when "1101110110100" => q_unbuf <= my_rom(7092);
      when "1101110110101" => q_unbuf <= my_rom(7093);
      when "1101110110110" => q_unbuf <= my_rom(7094);
      when "1101110110111" => q_unbuf <= my_rom(7095);
      when "1101110111000" => q_unbuf <= my_rom(7096);
      when "1101110111001" => q_unbuf <= my_rom(7097);
      when "1101110111010" => q_unbuf <= my_rom(7098);
      when "1101110111011" => q_unbuf <= my_rom(7099);
      when "1101110111100" => q_unbuf <= my_rom(7100);
      when "1101110111101" => q_unbuf <= my_rom(7101);
      when "1101110111110" => q_unbuf <= my_rom(7102);
      when "1101110111111" => q_unbuf <= my_rom(7103);
      when "1101111000000" => q_unbuf <= my_rom(7104);
      when "1101111000001" => q_unbuf <= my_rom(7105);
      when "1101111000010" => q_unbuf <= my_rom(7106);
      when "1101111000011" => q_unbuf <= my_rom(7107);
      when "1101111000100" => q_unbuf <= my_rom(7108);
      when "1101111000101" => q_unbuf <= my_rom(7109);
      when "1101111000110" => q_unbuf <= my_rom(7110);
      when "1101111000111" => q_unbuf <= my_rom(7111);
      when "1101111001000" => q_unbuf <= my_rom(7112);
      when "1101111001001" => q_unbuf <= my_rom(7113);
      when "1101111001010" => q_unbuf <= my_rom(7114);
      when "1101111001011" => q_unbuf <= my_rom(7115);
      when "1101111001100" => q_unbuf <= my_rom(7116);
      when "1101111001101" => q_unbuf <= my_rom(7117);
      when "1101111001110" => q_unbuf <= my_rom(7118);
      when "1101111001111" => q_unbuf <= my_rom(7119);
      when "1101111010000" => q_unbuf <= my_rom(7120);
      when "1101111010001" => q_unbuf <= my_rom(7121);
      when "1101111010010" => q_unbuf <= my_rom(7122);
      when "1101111010011" => q_unbuf <= my_rom(7123);
      when "1101111010100" => q_unbuf <= my_rom(7124);
      when "1101111010101" => q_unbuf <= my_rom(7125);
      when "1101111010110" => q_unbuf <= my_rom(7126);
      when "1101111010111" => q_unbuf <= my_rom(7127);
      when "1101111011000" => q_unbuf <= my_rom(7128);
      when "1101111011001" => q_unbuf <= my_rom(7129);
      when "1101111011010" => q_unbuf <= my_rom(7130);
      when "1101111011011" => q_unbuf <= my_rom(7131);
      when "1101111011100" => q_unbuf <= my_rom(7132);
      when "1101111011101" => q_unbuf <= my_rom(7133);
      when "1101111011110" => q_unbuf <= my_rom(7134);
      when "1101111011111" => q_unbuf <= my_rom(7135);
      when "1101111100000" => q_unbuf <= my_rom(7136);
      when "1101111100001" => q_unbuf <= my_rom(7137);
      when "1101111100010" => q_unbuf <= my_rom(7138);
      when "1101111100011" => q_unbuf <= my_rom(7139);
      when "1101111100100" => q_unbuf <= my_rom(7140);
      when "1101111100101" => q_unbuf <= my_rom(7141);
      when "1101111100110" => q_unbuf <= my_rom(7142);
      when "1101111100111" => q_unbuf <= my_rom(7143);
      when "1101111101000" => q_unbuf <= my_rom(7144);
      when "1101111101001" => q_unbuf <= my_rom(7145);
      when "1101111101010" => q_unbuf <= my_rom(7146);
      when "1101111101011" => q_unbuf <= my_rom(7147);
      when "1101111101100" => q_unbuf <= my_rom(7148);
      when "1101111101101" => q_unbuf <= my_rom(7149);
      when "1101111101110" => q_unbuf <= my_rom(7150);
      when "1101111101111" => q_unbuf <= my_rom(7151);
      when "1101111110000" => q_unbuf <= my_rom(7152);
      when "1101111110001" => q_unbuf <= my_rom(7153);
      when "1101111110010" => q_unbuf <= my_rom(7154);
      when "1101111110011" => q_unbuf <= my_rom(7155);
      when "1101111110100" => q_unbuf <= my_rom(7156);
      when "1101111110101" => q_unbuf <= my_rom(7157);
      when "1101111110110" => q_unbuf <= my_rom(7158);
      when "1101111110111" => q_unbuf <= my_rom(7159);
      when "1101111111000" => q_unbuf <= my_rom(7160);
      when "1101111111001" => q_unbuf <= my_rom(7161);
      when "1101111111010" => q_unbuf <= my_rom(7162);
      when "1101111111011" => q_unbuf <= my_rom(7163);
      when "1101111111100" => q_unbuf <= my_rom(7164);
      when "1101111111101" => q_unbuf <= my_rom(7165);
      when "1101111111110" => q_unbuf <= my_rom(7166);
      when "1101111111111" => q_unbuf <= my_rom(7167);
      when "1110000000000" => q_unbuf <= my_rom(7168);
      when "1110000000001" => q_unbuf <= my_rom(7169);
      when "1110000000010" => q_unbuf <= my_rom(7170);
      when "1110000000011" => q_unbuf <= my_rom(7171);
      when "1110000000100" => q_unbuf <= my_rom(7172);
      when "1110000000101" => q_unbuf <= my_rom(7173);
      when "1110000000110" => q_unbuf <= my_rom(7174);
      when "1110000000111" => q_unbuf <= my_rom(7175);
      when "1110000001000" => q_unbuf <= my_rom(7176);
      when "1110000001001" => q_unbuf <= my_rom(7177);
      when "1110000001010" => q_unbuf <= my_rom(7178);
      when "1110000001011" => q_unbuf <= my_rom(7179);
      when "1110000001100" => q_unbuf <= my_rom(7180);
      when "1110000001101" => q_unbuf <= my_rom(7181);
      when "1110000001110" => q_unbuf <= my_rom(7182);
      when "1110000001111" => q_unbuf <= my_rom(7183);
      when "1110000010000" => q_unbuf <= my_rom(7184);
      when "1110000010001" => q_unbuf <= my_rom(7185);
      when "1110000010010" => q_unbuf <= my_rom(7186);
      when "1110000010011" => q_unbuf <= my_rom(7187);
      when "1110000010100" => q_unbuf <= my_rom(7188);
      when "1110000010101" => q_unbuf <= my_rom(7189);
      when "1110000010110" => q_unbuf <= my_rom(7190);
      when "1110000010111" => q_unbuf <= my_rom(7191);
      when "1110000011000" => q_unbuf <= my_rom(7192);
      when "1110000011001" => q_unbuf <= my_rom(7193);
      when "1110000011010" => q_unbuf <= my_rom(7194);
      when "1110000011011" => q_unbuf <= my_rom(7195);
      when "1110000011100" => q_unbuf <= my_rom(7196);
      when "1110000011101" => q_unbuf <= my_rom(7197);
      when "1110000011110" => q_unbuf <= my_rom(7198);
      when "1110000011111" => q_unbuf <= my_rom(7199);
      when "1110000100000" => q_unbuf <= my_rom(7200);
      when "1110000100001" => q_unbuf <= my_rom(7201);
      when "1110000100010" => q_unbuf <= my_rom(7202);
      when "1110000100011" => q_unbuf <= my_rom(7203);
      when "1110000100100" => q_unbuf <= my_rom(7204);
      when "1110000100101" => q_unbuf <= my_rom(7205);
      when "1110000100110" => q_unbuf <= my_rom(7206);
      when "1110000100111" => q_unbuf <= my_rom(7207);
      when "1110000101000" => q_unbuf <= my_rom(7208);
      when "1110000101001" => q_unbuf <= my_rom(7209);
      when "1110000101010" => q_unbuf <= my_rom(7210);
      when "1110000101011" => q_unbuf <= my_rom(7211);
      when "1110000101100" => q_unbuf <= my_rom(7212);
      when "1110000101101" => q_unbuf <= my_rom(7213);
      when "1110000101110" => q_unbuf <= my_rom(7214);
      when "1110000101111" => q_unbuf <= my_rom(7215);
      when "1110000110000" => q_unbuf <= my_rom(7216);
      when "1110000110001" => q_unbuf <= my_rom(7217);
      when "1110000110010" => q_unbuf <= my_rom(7218);
      when "1110000110011" => q_unbuf <= my_rom(7219);
      when "1110000110100" => q_unbuf <= my_rom(7220);
      when "1110000110101" => q_unbuf <= my_rom(7221);
      when "1110000110110" => q_unbuf <= my_rom(7222);
      when "1110000110111" => q_unbuf <= my_rom(7223);
      when "1110000111000" => q_unbuf <= my_rom(7224);
      when "1110000111001" => q_unbuf <= my_rom(7225);
      when "1110000111010" => q_unbuf <= my_rom(7226);
      when "1110000111011" => q_unbuf <= my_rom(7227);
      when "1110000111100" => q_unbuf <= my_rom(7228);
      when "1110000111101" => q_unbuf <= my_rom(7229);
      when "1110000111110" => q_unbuf <= my_rom(7230);
      when "1110000111111" => q_unbuf <= my_rom(7231);
      when "1110001000000" => q_unbuf <= my_rom(7232);
      when "1110001000001" => q_unbuf <= my_rom(7233);
      when "1110001000010" => q_unbuf <= my_rom(7234);
      when "1110001000011" => q_unbuf <= my_rom(7235);
      when "1110001000100" => q_unbuf <= my_rom(7236);
      when "1110001000101" => q_unbuf <= my_rom(7237);
      when "1110001000110" => q_unbuf <= my_rom(7238);
      when "1110001000111" => q_unbuf <= my_rom(7239);
      when "1110001001000" => q_unbuf <= my_rom(7240);
      when "1110001001001" => q_unbuf <= my_rom(7241);
      when "1110001001010" => q_unbuf <= my_rom(7242);
      when "1110001001011" => q_unbuf <= my_rom(7243);
      when "1110001001100" => q_unbuf <= my_rom(7244);
      when "1110001001101" => q_unbuf <= my_rom(7245);
      when "1110001001110" => q_unbuf <= my_rom(7246);
      when "1110001001111" => q_unbuf <= my_rom(7247);
      when "1110001010000" => q_unbuf <= my_rom(7248);
      when "1110001010001" => q_unbuf <= my_rom(7249);
      when "1110001010010" => q_unbuf <= my_rom(7250);
      when "1110001010011" => q_unbuf <= my_rom(7251);
      when "1110001010100" => q_unbuf <= my_rom(7252);
      when "1110001010101" => q_unbuf <= my_rom(7253);
      when "1110001010110" => q_unbuf <= my_rom(7254);
      when "1110001010111" => q_unbuf <= my_rom(7255);
      when "1110001011000" => q_unbuf <= my_rom(7256);
      when "1110001011001" => q_unbuf <= my_rom(7257);
      when "1110001011010" => q_unbuf <= my_rom(7258);
      when "1110001011011" => q_unbuf <= my_rom(7259);
      when "1110001011100" => q_unbuf <= my_rom(7260);
      when "1110001011101" => q_unbuf <= my_rom(7261);
      when "1110001011110" => q_unbuf <= my_rom(7262);
      when "1110001011111" => q_unbuf <= my_rom(7263);
      when "1110001100000" => q_unbuf <= my_rom(7264);
      when "1110001100001" => q_unbuf <= my_rom(7265);
      when "1110001100010" => q_unbuf <= my_rom(7266);
      when "1110001100011" => q_unbuf <= my_rom(7267);
      when "1110001100100" => q_unbuf <= my_rom(7268);
      when "1110001100101" => q_unbuf <= my_rom(7269);
      when "1110001100110" => q_unbuf <= my_rom(7270);
      when "1110001100111" => q_unbuf <= my_rom(7271);
      when "1110001101000" => q_unbuf <= my_rom(7272);
      when "1110001101001" => q_unbuf <= my_rom(7273);
      when "1110001101010" => q_unbuf <= my_rom(7274);
      when "1110001101011" => q_unbuf <= my_rom(7275);
      when "1110001101100" => q_unbuf <= my_rom(7276);
      when "1110001101101" => q_unbuf <= my_rom(7277);
      when "1110001101110" => q_unbuf <= my_rom(7278);
      when "1110001101111" => q_unbuf <= my_rom(7279);
      when "1110001110000" => q_unbuf <= my_rom(7280);
      when "1110001110001" => q_unbuf <= my_rom(7281);
      when "1110001110010" => q_unbuf <= my_rom(7282);
      when "1110001110011" => q_unbuf <= my_rom(7283);
      when "1110001110100" => q_unbuf <= my_rom(7284);
      when "1110001110101" => q_unbuf <= my_rom(7285);
      when "1110001110110" => q_unbuf <= my_rom(7286);
      when "1110001110111" => q_unbuf <= my_rom(7287);
      when "1110001111000" => q_unbuf <= my_rom(7288);
      when "1110001111001" => q_unbuf <= my_rom(7289);
      when "1110001111010" => q_unbuf <= my_rom(7290);
      when "1110001111011" => q_unbuf <= my_rom(7291);
      when "1110001111100" => q_unbuf <= my_rom(7292);
      when "1110001111101" => q_unbuf <= my_rom(7293);
      when "1110001111110" => q_unbuf <= my_rom(7294);
      when "1110001111111" => q_unbuf <= my_rom(7295);
      when "1110010000000" => q_unbuf <= my_rom(7296);
      when "1110010000001" => q_unbuf <= my_rom(7297);
      when "1110010000010" => q_unbuf <= my_rom(7298);
      when "1110010000011" => q_unbuf <= my_rom(7299);
      when "1110010000100" => q_unbuf <= my_rom(7300);
      when "1110010000101" => q_unbuf <= my_rom(7301);
      when "1110010000110" => q_unbuf <= my_rom(7302);
      when "1110010000111" => q_unbuf <= my_rom(7303);
      when "1110010001000" => q_unbuf <= my_rom(7304);
      when "1110010001001" => q_unbuf <= my_rom(7305);
      when "1110010001010" => q_unbuf <= my_rom(7306);
      when "1110010001011" => q_unbuf <= my_rom(7307);
      when "1110010001100" => q_unbuf <= my_rom(7308);
      when "1110010001101" => q_unbuf <= my_rom(7309);
      when "1110010001110" => q_unbuf <= my_rom(7310);
      when "1110010001111" => q_unbuf <= my_rom(7311);
      when "1110010010000" => q_unbuf <= my_rom(7312);
      when "1110010010001" => q_unbuf <= my_rom(7313);
      when "1110010010010" => q_unbuf <= my_rom(7314);
      when "1110010010011" => q_unbuf <= my_rom(7315);
      when "1110010010100" => q_unbuf <= my_rom(7316);
      when "1110010010101" => q_unbuf <= my_rom(7317);
      when "1110010010110" => q_unbuf <= my_rom(7318);
      when "1110010010111" => q_unbuf <= my_rom(7319);
      when "1110010011000" => q_unbuf <= my_rom(7320);
      when "1110010011001" => q_unbuf <= my_rom(7321);
      when "1110010011010" => q_unbuf <= my_rom(7322);
      when "1110010011011" => q_unbuf <= my_rom(7323);
      when "1110010011100" => q_unbuf <= my_rom(7324);
      when "1110010011101" => q_unbuf <= my_rom(7325);
      when "1110010011110" => q_unbuf <= my_rom(7326);
      when "1110010011111" => q_unbuf <= my_rom(7327);
      when "1110010100000" => q_unbuf <= my_rom(7328);
      when "1110010100001" => q_unbuf <= my_rom(7329);
      when "1110010100010" => q_unbuf <= my_rom(7330);
      when "1110010100011" => q_unbuf <= my_rom(7331);
      when "1110010100100" => q_unbuf <= my_rom(7332);
      when "1110010100101" => q_unbuf <= my_rom(7333);
      when "1110010100110" => q_unbuf <= my_rom(7334);
      when "1110010100111" => q_unbuf <= my_rom(7335);
      when "1110010101000" => q_unbuf <= my_rom(7336);
      when "1110010101001" => q_unbuf <= my_rom(7337);
      when "1110010101010" => q_unbuf <= my_rom(7338);
      when "1110010101011" => q_unbuf <= my_rom(7339);
      when "1110010101100" => q_unbuf <= my_rom(7340);
      when "1110010101101" => q_unbuf <= my_rom(7341);
      when "1110010101110" => q_unbuf <= my_rom(7342);
      when "1110010101111" => q_unbuf <= my_rom(7343);
      when "1110010110000" => q_unbuf <= my_rom(7344);
      when "1110010110001" => q_unbuf <= my_rom(7345);
      when "1110010110010" => q_unbuf <= my_rom(7346);
      when "1110010110011" => q_unbuf <= my_rom(7347);
      when "1110010110100" => q_unbuf <= my_rom(7348);
      when "1110010110101" => q_unbuf <= my_rom(7349);
      when "1110010110110" => q_unbuf <= my_rom(7350);
      when "1110010110111" => q_unbuf <= my_rom(7351);
      when "1110010111000" => q_unbuf <= my_rom(7352);
      when "1110010111001" => q_unbuf <= my_rom(7353);
      when "1110010111010" => q_unbuf <= my_rom(7354);
      when "1110010111011" => q_unbuf <= my_rom(7355);
      when "1110010111100" => q_unbuf <= my_rom(7356);
      when "1110010111101" => q_unbuf <= my_rom(7357);
      when "1110010111110" => q_unbuf <= my_rom(7358);
      when "1110010111111" => q_unbuf <= my_rom(7359);
      when "1110011000000" => q_unbuf <= my_rom(7360);
      when "1110011000001" => q_unbuf <= my_rom(7361);
      when "1110011000010" => q_unbuf <= my_rom(7362);
      when "1110011000011" => q_unbuf <= my_rom(7363);
      when "1110011000100" => q_unbuf <= my_rom(7364);
      when "1110011000101" => q_unbuf <= my_rom(7365);
      when "1110011000110" => q_unbuf <= my_rom(7366);
      when "1110011000111" => q_unbuf <= my_rom(7367);
      when "1110011001000" => q_unbuf <= my_rom(7368);
      when "1110011001001" => q_unbuf <= my_rom(7369);
      when "1110011001010" => q_unbuf <= my_rom(7370);
      when "1110011001011" => q_unbuf <= my_rom(7371);
      when "1110011001100" => q_unbuf <= my_rom(7372);
      when "1110011001101" => q_unbuf <= my_rom(7373);
      when "1110011001110" => q_unbuf <= my_rom(7374);
      when "1110011001111" => q_unbuf <= my_rom(7375);
      when "1110011010000" => q_unbuf <= my_rom(7376);
      when "1110011010001" => q_unbuf <= my_rom(7377);
      when "1110011010010" => q_unbuf <= my_rom(7378);
      when "1110011010011" => q_unbuf <= my_rom(7379);
      when "1110011010100" => q_unbuf <= my_rom(7380);
      when "1110011010101" => q_unbuf <= my_rom(7381);
      when "1110011010110" => q_unbuf <= my_rom(7382);
      when "1110011010111" => q_unbuf <= my_rom(7383);
      when "1110011011000" => q_unbuf <= my_rom(7384);
      when "1110011011001" => q_unbuf <= my_rom(7385);
      when "1110011011010" => q_unbuf <= my_rom(7386);
      when "1110011011011" => q_unbuf <= my_rom(7387);
      when "1110011011100" => q_unbuf <= my_rom(7388);
      when "1110011011101" => q_unbuf <= my_rom(7389);
      when "1110011011110" => q_unbuf <= my_rom(7390);
      when "1110011011111" => q_unbuf <= my_rom(7391);
      when "1110011100000" => q_unbuf <= my_rom(7392);
      when "1110011100001" => q_unbuf <= my_rom(7393);
      when "1110011100010" => q_unbuf <= my_rom(7394);
      when "1110011100011" => q_unbuf <= my_rom(7395);
      when "1110011100100" => q_unbuf <= my_rom(7396);
      when "1110011100101" => q_unbuf <= my_rom(7397);
      when "1110011100110" => q_unbuf <= my_rom(7398);
      when "1110011100111" => q_unbuf <= my_rom(7399);
      when "1110011101000" => q_unbuf <= my_rom(7400);
      when "1110011101001" => q_unbuf <= my_rom(7401);
      when "1110011101010" => q_unbuf <= my_rom(7402);
      when "1110011101011" => q_unbuf <= my_rom(7403);
      when "1110011101100" => q_unbuf <= my_rom(7404);
      when "1110011101101" => q_unbuf <= my_rom(7405);
      when "1110011101110" => q_unbuf <= my_rom(7406);
      when "1110011101111" => q_unbuf <= my_rom(7407);
      when "1110011110000" => q_unbuf <= my_rom(7408);
      when "1110011110001" => q_unbuf <= my_rom(7409);
      when "1110011110010" => q_unbuf <= my_rom(7410);
      when "1110011110011" => q_unbuf <= my_rom(7411);
      when "1110011110100" => q_unbuf <= my_rom(7412);
      when "1110011110101" => q_unbuf <= my_rom(7413);
      when "1110011110110" => q_unbuf <= my_rom(7414);
      when "1110011110111" => q_unbuf <= my_rom(7415);
      when "1110011111000" => q_unbuf <= my_rom(7416);
      when "1110011111001" => q_unbuf <= my_rom(7417);
      when "1110011111010" => q_unbuf <= my_rom(7418);
      when "1110011111011" => q_unbuf <= my_rom(7419);
      when "1110011111100" => q_unbuf <= my_rom(7420);
      when "1110011111101" => q_unbuf <= my_rom(7421);
      when "1110011111110" => q_unbuf <= my_rom(7422);
      when "1110011111111" => q_unbuf <= my_rom(7423);
      when "1110100000000" => q_unbuf <= my_rom(7424);
      when "1110100000001" => q_unbuf <= my_rom(7425);
      when "1110100000010" => q_unbuf <= my_rom(7426);
      when "1110100000011" => q_unbuf <= my_rom(7427);
      when "1110100000100" => q_unbuf <= my_rom(7428);
      when "1110100000101" => q_unbuf <= my_rom(7429);
      when "1110100000110" => q_unbuf <= my_rom(7430);
      when "1110100000111" => q_unbuf <= my_rom(7431);
      when "1110100001000" => q_unbuf <= my_rom(7432);
      when "1110100001001" => q_unbuf <= my_rom(7433);
      when "1110100001010" => q_unbuf <= my_rom(7434);
      when "1110100001011" => q_unbuf <= my_rom(7435);
      when "1110100001100" => q_unbuf <= my_rom(7436);
      when "1110100001101" => q_unbuf <= my_rom(7437);
      when "1110100001110" => q_unbuf <= my_rom(7438);
      when "1110100001111" => q_unbuf <= my_rom(7439);
      when "1110100010000" => q_unbuf <= my_rom(7440);
      when "1110100010001" => q_unbuf <= my_rom(7441);
      when "1110100010010" => q_unbuf <= my_rom(7442);
      when "1110100010011" => q_unbuf <= my_rom(7443);
      when "1110100010100" => q_unbuf <= my_rom(7444);
      when "1110100010101" => q_unbuf <= my_rom(7445);
      when "1110100010110" => q_unbuf <= my_rom(7446);
      when "1110100010111" => q_unbuf <= my_rom(7447);
      when "1110100011000" => q_unbuf <= my_rom(7448);
      when "1110100011001" => q_unbuf <= my_rom(7449);
      when "1110100011010" => q_unbuf <= my_rom(7450);
      when "1110100011011" => q_unbuf <= my_rom(7451);
      when "1110100011100" => q_unbuf <= my_rom(7452);
      when "1110100011101" => q_unbuf <= my_rom(7453);
      when "1110100011110" => q_unbuf <= my_rom(7454);
      when "1110100011111" => q_unbuf <= my_rom(7455);
      when "1110100100000" => q_unbuf <= my_rom(7456);
      when "1110100100001" => q_unbuf <= my_rom(7457);
      when "1110100100010" => q_unbuf <= my_rom(7458);
      when "1110100100011" => q_unbuf <= my_rom(7459);
      when "1110100100100" => q_unbuf <= my_rom(7460);
      when "1110100100101" => q_unbuf <= my_rom(7461);
      when "1110100100110" => q_unbuf <= my_rom(7462);
      when "1110100100111" => q_unbuf <= my_rom(7463);
      when "1110100101000" => q_unbuf <= my_rom(7464);
      when "1110100101001" => q_unbuf <= my_rom(7465);
      when "1110100101010" => q_unbuf <= my_rom(7466);
      when "1110100101011" => q_unbuf <= my_rom(7467);
      when "1110100101100" => q_unbuf <= my_rom(7468);
      when "1110100101101" => q_unbuf <= my_rom(7469);
      when "1110100101110" => q_unbuf <= my_rom(7470);
      when "1110100101111" => q_unbuf <= my_rom(7471);
      when "1110100110000" => q_unbuf <= my_rom(7472);
      when "1110100110001" => q_unbuf <= my_rom(7473);
      when "1110100110010" => q_unbuf <= my_rom(7474);
      when "1110100110011" => q_unbuf <= my_rom(7475);
      when "1110100110100" => q_unbuf <= my_rom(7476);
      when "1110100110101" => q_unbuf <= my_rom(7477);
      when "1110100110110" => q_unbuf <= my_rom(7478);
      when "1110100110111" => q_unbuf <= my_rom(7479);
      when "1110100111000" => q_unbuf <= my_rom(7480);
      when "1110100111001" => q_unbuf <= my_rom(7481);
      when "1110100111010" => q_unbuf <= my_rom(7482);
      when "1110100111011" => q_unbuf <= my_rom(7483);
      when "1110100111100" => q_unbuf <= my_rom(7484);
      when "1110100111101" => q_unbuf <= my_rom(7485);
      when "1110100111110" => q_unbuf <= my_rom(7486);
      when "1110100111111" => q_unbuf <= my_rom(7487);
      when "1110101000000" => q_unbuf <= my_rom(7488);
      when "1110101000001" => q_unbuf <= my_rom(7489);
      when "1110101000010" => q_unbuf <= my_rom(7490);
      when "1110101000011" => q_unbuf <= my_rom(7491);
      when "1110101000100" => q_unbuf <= my_rom(7492);
      when "1110101000101" => q_unbuf <= my_rom(7493);
      when "1110101000110" => q_unbuf <= my_rom(7494);
      when "1110101000111" => q_unbuf <= my_rom(7495);
      when "1110101001000" => q_unbuf <= my_rom(7496);
      when "1110101001001" => q_unbuf <= my_rom(7497);
      when "1110101001010" => q_unbuf <= my_rom(7498);
      when "1110101001011" => q_unbuf <= my_rom(7499);
      when "1110101001100" => q_unbuf <= my_rom(7500);
      when "1110101001101" => q_unbuf <= my_rom(7501);
      when "1110101001110" => q_unbuf <= my_rom(7502);
      when "1110101001111" => q_unbuf <= my_rom(7503);
      when "1110101010000" => q_unbuf <= my_rom(7504);
      when "1110101010001" => q_unbuf <= my_rom(7505);
      when "1110101010010" => q_unbuf <= my_rom(7506);
      when "1110101010011" => q_unbuf <= my_rom(7507);
      when "1110101010100" => q_unbuf <= my_rom(7508);
      when "1110101010101" => q_unbuf <= my_rom(7509);
      when "1110101010110" => q_unbuf <= my_rom(7510);
      when "1110101010111" => q_unbuf <= my_rom(7511);
      when "1110101011000" => q_unbuf <= my_rom(7512);
      when "1110101011001" => q_unbuf <= my_rom(7513);
      when "1110101011010" => q_unbuf <= my_rom(7514);
      when "1110101011011" => q_unbuf <= my_rom(7515);
      when "1110101011100" => q_unbuf <= my_rom(7516);
      when "1110101011101" => q_unbuf <= my_rom(7517);
      when "1110101011110" => q_unbuf <= my_rom(7518);
      when "1110101011111" => q_unbuf <= my_rom(7519);
      when "1110101100000" => q_unbuf <= my_rom(7520);
      when "1110101100001" => q_unbuf <= my_rom(7521);
      when "1110101100010" => q_unbuf <= my_rom(7522);
      when "1110101100011" => q_unbuf <= my_rom(7523);
      when "1110101100100" => q_unbuf <= my_rom(7524);
      when "1110101100101" => q_unbuf <= my_rom(7525);
      when "1110101100110" => q_unbuf <= my_rom(7526);
      when "1110101100111" => q_unbuf <= my_rom(7527);
      when "1110101101000" => q_unbuf <= my_rom(7528);
      when "1110101101001" => q_unbuf <= my_rom(7529);
      when "1110101101010" => q_unbuf <= my_rom(7530);
      when "1110101101011" => q_unbuf <= my_rom(7531);
      when "1110101101100" => q_unbuf <= my_rom(7532);
      when "1110101101101" => q_unbuf <= my_rom(7533);
      when "1110101101110" => q_unbuf <= my_rom(7534);
      when "1110101101111" => q_unbuf <= my_rom(7535);
      when "1110101110000" => q_unbuf <= my_rom(7536);
      when "1110101110001" => q_unbuf <= my_rom(7537);
      when "1110101110010" => q_unbuf <= my_rom(7538);
      when "1110101110011" => q_unbuf <= my_rom(7539);
      when "1110101110100" => q_unbuf <= my_rom(7540);
      when "1110101110101" => q_unbuf <= my_rom(7541);
      when "1110101110110" => q_unbuf <= my_rom(7542);
      when "1110101110111" => q_unbuf <= my_rom(7543);
      when "1110101111000" => q_unbuf <= my_rom(7544);
      when "1110101111001" => q_unbuf <= my_rom(7545);
      when "1110101111010" => q_unbuf <= my_rom(7546);
      when "1110101111011" => q_unbuf <= my_rom(7547);
      when "1110101111100" => q_unbuf <= my_rom(7548);
      when "1110101111101" => q_unbuf <= my_rom(7549);
      when "1110101111110" => q_unbuf <= my_rom(7550);
      when "1110101111111" => q_unbuf <= my_rom(7551);
      when "1110110000000" => q_unbuf <= my_rom(7552);
      when "1110110000001" => q_unbuf <= my_rom(7553);
      when "1110110000010" => q_unbuf <= my_rom(7554);
      when "1110110000011" => q_unbuf <= my_rom(7555);
      when "1110110000100" => q_unbuf <= my_rom(7556);
      when "1110110000101" => q_unbuf <= my_rom(7557);
      when "1110110000110" => q_unbuf <= my_rom(7558);
      when "1110110000111" => q_unbuf <= my_rom(7559);
      when "1110110001000" => q_unbuf <= my_rom(7560);
      when "1110110001001" => q_unbuf <= my_rom(7561);
      when "1110110001010" => q_unbuf <= my_rom(7562);
      when "1110110001011" => q_unbuf <= my_rom(7563);
      when "1110110001100" => q_unbuf <= my_rom(7564);
      when "1110110001101" => q_unbuf <= my_rom(7565);
      when "1110110001110" => q_unbuf <= my_rom(7566);
      when "1110110001111" => q_unbuf <= my_rom(7567);
      when "1110110010000" => q_unbuf <= my_rom(7568);
      when "1110110010001" => q_unbuf <= my_rom(7569);
      when "1110110010010" => q_unbuf <= my_rom(7570);
      when "1110110010011" => q_unbuf <= my_rom(7571);
      when "1110110010100" => q_unbuf <= my_rom(7572);
      when "1110110010101" => q_unbuf <= my_rom(7573);
      when "1110110010110" => q_unbuf <= my_rom(7574);
      when "1110110010111" => q_unbuf <= my_rom(7575);
      when "1110110011000" => q_unbuf <= my_rom(7576);
      when "1110110011001" => q_unbuf <= my_rom(7577);
      when "1110110011010" => q_unbuf <= my_rom(7578);
      when "1110110011011" => q_unbuf <= my_rom(7579);
      when "1110110011100" => q_unbuf <= my_rom(7580);
      when "1110110011101" => q_unbuf <= my_rom(7581);
      when "1110110011110" => q_unbuf <= my_rom(7582);
      when "1110110011111" => q_unbuf <= my_rom(7583);
      when "1110110100000" => q_unbuf <= my_rom(7584);
      when "1110110100001" => q_unbuf <= my_rom(7585);
      when "1110110100010" => q_unbuf <= my_rom(7586);
      when "1110110100011" => q_unbuf <= my_rom(7587);
      when "1110110100100" => q_unbuf <= my_rom(7588);
      when "1110110100101" => q_unbuf <= my_rom(7589);
      when "1110110100110" => q_unbuf <= my_rom(7590);
      when "1110110100111" => q_unbuf <= my_rom(7591);
      when "1110110101000" => q_unbuf <= my_rom(7592);
      when "1110110101001" => q_unbuf <= my_rom(7593);
      when "1110110101010" => q_unbuf <= my_rom(7594);
      when "1110110101011" => q_unbuf <= my_rom(7595);
      when "1110110101100" => q_unbuf <= my_rom(7596);
      when "1110110101101" => q_unbuf <= my_rom(7597);
      when "1110110101110" => q_unbuf <= my_rom(7598);
      when "1110110101111" => q_unbuf <= my_rom(7599);
      when "1110110110000" => q_unbuf <= my_rom(7600);
      when "1110110110001" => q_unbuf <= my_rom(7601);
      when "1110110110010" => q_unbuf <= my_rom(7602);
      when "1110110110011" => q_unbuf <= my_rom(7603);
      when "1110110110100" => q_unbuf <= my_rom(7604);
      when "1110110110101" => q_unbuf <= my_rom(7605);
      when "1110110110110" => q_unbuf <= my_rom(7606);
      when "1110110110111" => q_unbuf <= my_rom(7607);
      when "1110110111000" => q_unbuf <= my_rom(7608);
      when "1110110111001" => q_unbuf <= my_rom(7609);
      when "1110110111010" => q_unbuf <= my_rom(7610);
      when "1110110111011" => q_unbuf <= my_rom(7611);
      when "1110110111100" => q_unbuf <= my_rom(7612);
      when "1110110111101" => q_unbuf <= my_rom(7613);
      when "1110110111110" => q_unbuf <= my_rom(7614);
      when "1110110111111" => q_unbuf <= my_rom(7615);
      when "1110111000000" => q_unbuf <= my_rom(7616);
      when "1110111000001" => q_unbuf <= my_rom(7617);
      when "1110111000010" => q_unbuf <= my_rom(7618);
      when "1110111000011" => q_unbuf <= my_rom(7619);
      when "1110111000100" => q_unbuf <= my_rom(7620);
      when "1110111000101" => q_unbuf <= my_rom(7621);
      when "1110111000110" => q_unbuf <= my_rom(7622);
      when "1110111000111" => q_unbuf <= my_rom(7623);
      when "1110111001000" => q_unbuf <= my_rom(7624);
      when "1110111001001" => q_unbuf <= my_rom(7625);
      when "1110111001010" => q_unbuf <= my_rom(7626);
      when "1110111001011" => q_unbuf <= my_rom(7627);
      when "1110111001100" => q_unbuf <= my_rom(7628);
      when "1110111001101" => q_unbuf <= my_rom(7629);
      when "1110111001110" => q_unbuf <= my_rom(7630);
      when "1110111001111" => q_unbuf <= my_rom(7631);
      when "1110111010000" => q_unbuf <= my_rom(7632);
      when "1110111010001" => q_unbuf <= my_rom(7633);
      when "1110111010010" => q_unbuf <= my_rom(7634);
      when "1110111010011" => q_unbuf <= my_rom(7635);
      when "1110111010100" => q_unbuf <= my_rom(7636);
      when "1110111010101" => q_unbuf <= my_rom(7637);
      when "1110111010110" => q_unbuf <= my_rom(7638);
      when "1110111010111" => q_unbuf <= my_rom(7639);
      when "1110111011000" => q_unbuf <= my_rom(7640);
      when "1110111011001" => q_unbuf <= my_rom(7641);
      when "1110111011010" => q_unbuf <= my_rom(7642);
      when "1110111011011" => q_unbuf <= my_rom(7643);
      when "1110111011100" => q_unbuf <= my_rom(7644);
      when "1110111011101" => q_unbuf <= my_rom(7645);
      when "1110111011110" => q_unbuf <= my_rom(7646);
      when "1110111011111" => q_unbuf <= my_rom(7647);
      when "1110111100000" => q_unbuf <= my_rom(7648);
      when "1110111100001" => q_unbuf <= my_rom(7649);
      when "1110111100010" => q_unbuf <= my_rom(7650);
      when "1110111100011" => q_unbuf <= my_rom(7651);
      when "1110111100100" => q_unbuf <= my_rom(7652);
      when "1110111100101" => q_unbuf <= my_rom(7653);
      when "1110111100110" => q_unbuf <= my_rom(7654);
      when "1110111100111" => q_unbuf <= my_rom(7655);
      when "1110111101000" => q_unbuf <= my_rom(7656);
      when "1110111101001" => q_unbuf <= my_rom(7657);
      when "1110111101010" => q_unbuf <= my_rom(7658);
      when "1110111101011" => q_unbuf <= my_rom(7659);
      when "1110111101100" => q_unbuf <= my_rom(7660);
      when "1110111101101" => q_unbuf <= my_rom(7661);
      when "1110111101110" => q_unbuf <= my_rom(7662);
      when "1110111101111" => q_unbuf <= my_rom(7663);
      when "1110111110000" => q_unbuf <= my_rom(7664);
      when "1110111110001" => q_unbuf <= my_rom(7665);
      when "1110111110010" => q_unbuf <= my_rom(7666);
      when "1110111110011" => q_unbuf <= my_rom(7667);
      when "1110111110100" => q_unbuf <= my_rom(7668);
      when "1110111110101" => q_unbuf <= my_rom(7669);
      when "1110111110110" => q_unbuf <= my_rom(7670);
      when "1110111110111" => q_unbuf <= my_rom(7671);
      when "1110111111000" => q_unbuf <= my_rom(7672);
      when "1110111111001" => q_unbuf <= my_rom(7673);
      when "1110111111010" => q_unbuf <= my_rom(7674);
      when "1110111111011" => q_unbuf <= my_rom(7675);
      when "1110111111100" => q_unbuf <= my_rom(7676);
      when "1110111111101" => q_unbuf <= my_rom(7677);
      when "1110111111110" => q_unbuf <= my_rom(7678);
      when "1110111111111" => q_unbuf <= my_rom(7679);
      when "1111000000000" => q_unbuf <= my_rom(7680);
      when "1111000000001" => q_unbuf <= my_rom(7681);
      when "1111000000010" => q_unbuf <= my_rom(7682);
      when "1111000000011" => q_unbuf <= my_rom(7683);
      when "1111000000100" => q_unbuf <= my_rom(7684);
      when "1111000000101" => q_unbuf <= my_rom(7685);
      when "1111000000110" => q_unbuf <= my_rom(7686);
      when "1111000000111" => q_unbuf <= my_rom(7687);
      when "1111000001000" => q_unbuf <= my_rom(7688);
      when "1111000001001" => q_unbuf <= my_rom(7689);
      when "1111000001010" => q_unbuf <= my_rom(7690);
      when "1111000001011" => q_unbuf <= my_rom(7691);
      when "1111000001100" => q_unbuf <= my_rom(7692);
      when "1111000001101" => q_unbuf <= my_rom(7693);
      when "1111000001110" => q_unbuf <= my_rom(7694);
      when "1111000001111" => q_unbuf <= my_rom(7695);
      when "1111000010000" => q_unbuf <= my_rom(7696);
      when "1111000010001" => q_unbuf <= my_rom(7697);
      when "1111000010010" => q_unbuf <= my_rom(7698);
      when "1111000010011" => q_unbuf <= my_rom(7699);
      when "1111000010100" => q_unbuf <= my_rom(7700);
      when "1111000010101" => q_unbuf <= my_rom(7701);
      when "1111000010110" => q_unbuf <= my_rom(7702);
      when "1111000010111" => q_unbuf <= my_rom(7703);
      when "1111000011000" => q_unbuf <= my_rom(7704);
      when "1111000011001" => q_unbuf <= my_rom(7705);
      when "1111000011010" => q_unbuf <= my_rom(7706);
      when "1111000011011" => q_unbuf <= my_rom(7707);
      when "1111000011100" => q_unbuf <= my_rom(7708);
      when "1111000011101" => q_unbuf <= my_rom(7709);
      when "1111000011110" => q_unbuf <= my_rom(7710);
      when "1111000011111" => q_unbuf <= my_rom(7711);
      when "1111000100000" => q_unbuf <= my_rom(7712);
      when "1111000100001" => q_unbuf <= my_rom(7713);
      when "1111000100010" => q_unbuf <= my_rom(7714);
      when "1111000100011" => q_unbuf <= my_rom(7715);
      when "1111000100100" => q_unbuf <= my_rom(7716);
      when "1111000100101" => q_unbuf <= my_rom(7717);
      when "1111000100110" => q_unbuf <= my_rom(7718);
      when "1111000100111" => q_unbuf <= my_rom(7719);
      when "1111000101000" => q_unbuf <= my_rom(7720);
      when "1111000101001" => q_unbuf <= my_rom(7721);
      when "1111000101010" => q_unbuf <= my_rom(7722);
      when "1111000101011" => q_unbuf <= my_rom(7723);
      when "1111000101100" => q_unbuf <= my_rom(7724);
      when "1111000101101" => q_unbuf <= my_rom(7725);
      when "1111000101110" => q_unbuf <= my_rom(7726);
      when "1111000101111" => q_unbuf <= my_rom(7727);
      when "1111000110000" => q_unbuf <= my_rom(7728);
      when "1111000110001" => q_unbuf <= my_rom(7729);
      when "1111000110010" => q_unbuf <= my_rom(7730);
      when "1111000110011" => q_unbuf <= my_rom(7731);
      when "1111000110100" => q_unbuf <= my_rom(7732);
      when "1111000110101" => q_unbuf <= my_rom(7733);
      when "1111000110110" => q_unbuf <= my_rom(7734);
      when "1111000110111" => q_unbuf <= my_rom(7735);
      when "1111000111000" => q_unbuf <= my_rom(7736);
      when "1111000111001" => q_unbuf <= my_rom(7737);
      when "1111000111010" => q_unbuf <= my_rom(7738);
      when "1111000111011" => q_unbuf <= my_rom(7739);
      when "1111000111100" => q_unbuf <= my_rom(7740);
      when "1111000111101" => q_unbuf <= my_rom(7741);
      when "1111000111110" => q_unbuf <= my_rom(7742);
      when "1111000111111" => q_unbuf <= my_rom(7743);
      when "1111001000000" => q_unbuf <= my_rom(7744);
      when "1111001000001" => q_unbuf <= my_rom(7745);
      when "1111001000010" => q_unbuf <= my_rom(7746);
      when "1111001000011" => q_unbuf <= my_rom(7747);
      when "1111001000100" => q_unbuf <= my_rom(7748);
      when "1111001000101" => q_unbuf <= my_rom(7749);
      when "1111001000110" => q_unbuf <= my_rom(7750);
      when "1111001000111" => q_unbuf <= my_rom(7751);
      when "1111001001000" => q_unbuf <= my_rom(7752);
      when "1111001001001" => q_unbuf <= my_rom(7753);
      when "1111001001010" => q_unbuf <= my_rom(7754);
      when "1111001001011" => q_unbuf <= my_rom(7755);
      when "1111001001100" => q_unbuf <= my_rom(7756);
      when "1111001001101" => q_unbuf <= my_rom(7757);
      when "1111001001110" => q_unbuf <= my_rom(7758);
      when "1111001001111" => q_unbuf <= my_rom(7759);
      when "1111001010000" => q_unbuf <= my_rom(7760);
      when "1111001010001" => q_unbuf <= my_rom(7761);
      when "1111001010010" => q_unbuf <= my_rom(7762);
      when "1111001010011" => q_unbuf <= my_rom(7763);
      when "1111001010100" => q_unbuf <= my_rom(7764);
      when "1111001010101" => q_unbuf <= my_rom(7765);
      when "1111001010110" => q_unbuf <= my_rom(7766);
      when "1111001010111" => q_unbuf <= my_rom(7767);
      when "1111001011000" => q_unbuf <= my_rom(7768);
      when "1111001011001" => q_unbuf <= my_rom(7769);
      when "1111001011010" => q_unbuf <= my_rom(7770);
      when "1111001011011" => q_unbuf <= my_rom(7771);
      when "1111001011100" => q_unbuf <= my_rom(7772);
      when "1111001011101" => q_unbuf <= my_rom(7773);
      when "1111001011110" => q_unbuf <= my_rom(7774);
      when "1111001011111" => q_unbuf <= my_rom(7775);
      when "1111001100000" => q_unbuf <= my_rom(7776);
      when "1111001100001" => q_unbuf <= my_rom(7777);
      when "1111001100010" => q_unbuf <= my_rom(7778);
      when "1111001100011" => q_unbuf <= my_rom(7779);
      when "1111001100100" => q_unbuf <= my_rom(7780);
      when "1111001100101" => q_unbuf <= my_rom(7781);
      when "1111001100110" => q_unbuf <= my_rom(7782);
      when "1111001100111" => q_unbuf <= my_rom(7783);
      when "1111001101000" => q_unbuf <= my_rom(7784);
      when "1111001101001" => q_unbuf <= my_rom(7785);
      when "1111001101010" => q_unbuf <= my_rom(7786);
      when "1111001101011" => q_unbuf <= my_rom(7787);
      when "1111001101100" => q_unbuf <= my_rom(7788);
      when "1111001101101" => q_unbuf <= my_rom(7789);
      when "1111001101110" => q_unbuf <= my_rom(7790);
      when "1111001101111" => q_unbuf <= my_rom(7791);
      when "1111001110000" => q_unbuf <= my_rom(7792);
      when "1111001110001" => q_unbuf <= my_rom(7793);
      when "1111001110010" => q_unbuf <= my_rom(7794);
      when "1111001110011" => q_unbuf <= my_rom(7795);
      when "1111001110100" => q_unbuf <= my_rom(7796);
      when "1111001110101" => q_unbuf <= my_rom(7797);
      when "1111001110110" => q_unbuf <= my_rom(7798);
      when "1111001110111" => q_unbuf <= my_rom(7799);
      when "1111001111000" => q_unbuf <= my_rom(7800);
      when "1111001111001" => q_unbuf <= my_rom(7801);
      when "1111001111010" => q_unbuf <= my_rom(7802);
      when "1111001111011" => q_unbuf <= my_rom(7803);
      when "1111001111100" => q_unbuf <= my_rom(7804);
      when "1111001111101" => q_unbuf <= my_rom(7805);
      when "1111001111110" => q_unbuf <= my_rom(7806);
      when "1111001111111" => q_unbuf <= my_rom(7807);
      when "1111010000000" => q_unbuf <= my_rom(7808);
      when "1111010000001" => q_unbuf <= my_rom(7809);
      when "1111010000010" => q_unbuf <= my_rom(7810);
      when "1111010000011" => q_unbuf <= my_rom(7811);
      when "1111010000100" => q_unbuf <= my_rom(7812);
      when "1111010000101" => q_unbuf <= my_rom(7813);
      when "1111010000110" => q_unbuf <= my_rom(7814);
      when "1111010000111" => q_unbuf <= my_rom(7815);
      when "1111010001000" => q_unbuf <= my_rom(7816);
      when "1111010001001" => q_unbuf <= my_rom(7817);
      when "1111010001010" => q_unbuf <= my_rom(7818);
      when "1111010001011" => q_unbuf <= my_rom(7819);
      when "1111010001100" => q_unbuf <= my_rom(7820);
      when "1111010001101" => q_unbuf <= my_rom(7821);
      when "1111010001110" => q_unbuf <= my_rom(7822);
      when "1111010001111" => q_unbuf <= my_rom(7823);
      when "1111010010000" => q_unbuf <= my_rom(7824);
      when "1111010010001" => q_unbuf <= my_rom(7825);
      when "1111010010010" => q_unbuf <= my_rom(7826);
      when "1111010010011" => q_unbuf <= my_rom(7827);
      when "1111010010100" => q_unbuf <= my_rom(7828);
      when "1111010010101" => q_unbuf <= my_rom(7829);
      when "1111010010110" => q_unbuf <= my_rom(7830);
      when "1111010010111" => q_unbuf <= my_rom(7831);
      when "1111010011000" => q_unbuf <= my_rom(7832);
      when "1111010011001" => q_unbuf <= my_rom(7833);
      when "1111010011010" => q_unbuf <= my_rom(7834);
      when "1111010011011" => q_unbuf <= my_rom(7835);
      when "1111010011100" => q_unbuf <= my_rom(7836);
      when "1111010011101" => q_unbuf <= my_rom(7837);
      when "1111010011110" => q_unbuf <= my_rom(7838);
      when "1111010011111" => q_unbuf <= my_rom(7839);
      when "1111010100000" => q_unbuf <= my_rom(7840);
      when "1111010100001" => q_unbuf <= my_rom(7841);
      when "1111010100010" => q_unbuf <= my_rom(7842);
      when "1111010100011" => q_unbuf <= my_rom(7843);
      when "1111010100100" => q_unbuf <= my_rom(7844);
      when "1111010100101" => q_unbuf <= my_rom(7845);
      when "1111010100110" => q_unbuf <= my_rom(7846);
      when "1111010100111" => q_unbuf <= my_rom(7847);
      when "1111010101000" => q_unbuf <= my_rom(7848);
      when "1111010101001" => q_unbuf <= my_rom(7849);
      when "1111010101010" => q_unbuf <= my_rom(7850);
      when "1111010101011" => q_unbuf <= my_rom(7851);
      when "1111010101100" => q_unbuf <= my_rom(7852);
      when "1111010101101" => q_unbuf <= my_rom(7853);
      when "1111010101110" => q_unbuf <= my_rom(7854);
      when "1111010101111" => q_unbuf <= my_rom(7855);
      when "1111010110000" => q_unbuf <= my_rom(7856);
      when "1111010110001" => q_unbuf <= my_rom(7857);
      when "1111010110010" => q_unbuf <= my_rom(7858);
      when "1111010110011" => q_unbuf <= my_rom(7859);
      when "1111010110100" => q_unbuf <= my_rom(7860);
      when "1111010110101" => q_unbuf <= my_rom(7861);
      when "1111010110110" => q_unbuf <= my_rom(7862);
      when "1111010110111" => q_unbuf <= my_rom(7863);
      when "1111010111000" => q_unbuf <= my_rom(7864);
      when "1111010111001" => q_unbuf <= my_rom(7865);
      when "1111010111010" => q_unbuf <= my_rom(7866);
      when "1111010111011" => q_unbuf <= my_rom(7867);
      when "1111010111100" => q_unbuf <= my_rom(7868);
      when "1111010111101" => q_unbuf <= my_rom(7869);
      when "1111010111110" => q_unbuf <= my_rom(7870);
      when "1111010111111" => q_unbuf <= my_rom(7871);
      when "1111011000000" => q_unbuf <= my_rom(7872);
      when "1111011000001" => q_unbuf <= my_rom(7873);
      when "1111011000010" => q_unbuf <= my_rom(7874);
      when "1111011000011" => q_unbuf <= my_rom(7875);
      when "1111011000100" => q_unbuf <= my_rom(7876);
      when "1111011000101" => q_unbuf <= my_rom(7877);
      when "1111011000110" => q_unbuf <= my_rom(7878);
      when "1111011000111" => q_unbuf <= my_rom(7879);
      when "1111011001000" => q_unbuf <= my_rom(7880);
      when "1111011001001" => q_unbuf <= my_rom(7881);
      when "1111011001010" => q_unbuf <= my_rom(7882);
      when "1111011001011" => q_unbuf <= my_rom(7883);
      when "1111011001100" => q_unbuf <= my_rom(7884);
      when "1111011001101" => q_unbuf <= my_rom(7885);
      when "1111011001110" => q_unbuf <= my_rom(7886);
      when "1111011001111" => q_unbuf <= my_rom(7887);
      when "1111011010000" => q_unbuf <= my_rom(7888);
      when "1111011010001" => q_unbuf <= my_rom(7889);
      when "1111011010010" => q_unbuf <= my_rom(7890);
      when "1111011010011" => q_unbuf <= my_rom(7891);
      when "1111011010100" => q_unbuf <= my_rom(7892);
      when "1111011010101" => q_unbuf <= my_rom(7893);
      when "1111011010110" => q_unbuf <= my_rom(7894);
      when "1111011010111" => q_unbuf <= my_rom(7895);
      when "1111011011000" => q_unbuf <= my_rom(7896);
      when "1111011011001" => q_unbuf <= my_rom(7897);
      when "1111011011010" => q_unbuf <= my_rom(7898);
      when "1111011011011" => q_unbuf <= my_rom(7899);
      when "1111011011100" => q_unbuf <= my_rom(7900);
      when "1111011011101" => q_unbuf <= my_rom(7901);
      when "1111011011110" => q_unbuf <= my_rom(7902);
      when "1111011011111" => q_unbuf <= my_rom(7903);
      when "1111011100000" => q_unbuf <= my_rom(7904);
      when "1111011100001" => q_unbuf <= my_rom(7905);
      when "1111011100010" => q_unbuf <= my_rom(7906);
      when "1111011100011" => q_unbuf <= my_rom(7907);
      when "1111011100100" => q_unbuf <= my_rom(7908);
      when "1111011100101" => q_unbuf <= my_rom(7909);
      when "1111011100110" => q_unbuf <= my_rom(7910);
      when "1111011100111" => q_unbuf <= my_rom(7911);
      when "1111011101000" => q_unbuf <= my_rom(7912);
      when "1111011101001" => q_unbuf <= my_rom(7913);
      when "1111011101010" => q_unbuf <= my_rom(7914);
      when "1111011101011" => q_unbuf <= my_rom(7915);
      when "1111011101100" => q_unbuf <= my_rom(7916);
      when "1111011101101" => q_unbuf <= my_rom(7917);
      when "1111011101110" => q_unbuf <= my_rom(7918);
      when "1111011101111" => q_unbuf <= my_rom(7919);
      when "1111011110000" => q_unbuf <= my_rom(7920);
      when "1111011110001" => q_unbuf <= my_rom(7921);
      when "1111011110010" => q_unbuf <= my_rom(7922);
      when "1111011110011" => q_unbuf <= my_rom(7923);
      when "1111011110100" => q_unbuf <= my_rom(7924);
      when "1111011110101" => q_unbuf <= my_rom(7925);
      when "1111011110110" => q_unbuf <= my_rom(7926);
      when "1111011110111" => q_unbuf <= my_rom(7927);
      when "1111011111000" => q_unbuf <= my_rom(7928);
      when "1111011111001" => q_unbuf <= my_rom(7929);
      when "1111011111010" => q_unbuf <= my_rom(7930);
      when "1111011111011" => q_unbuf <= my_rom(7931);
      when "1111011111100" => q_unbuf <= my_rom(7932);
      when "1111011111101" => q_unbuf <= my_rom(7933);
      when "1111011111110" => q_unbuf <= my_rom(7934);
      when "1111011111111" => q_unbuf <= my_rom(7935);
      when "1111100000000" => q_unbuf <= my_rom(7936);
      when "1111100000001" => q_unbuf <= my_rom(7937);
      when "1111100000010" => q_unbuf <= my_rom(7938);
      when "1111100000011" => q_unbuf <= my_rom(7939);
      when "1111100000100" => q_unbuf <= my_rom(7940);
      when "1111100000101" => q_unbuf <= my_rom(7941);
      when "1111100000110" => q_unbuf <= my_rom(7942);
      when "1111100000111" => q_unbuf <= my_rom(7943);
      when "1111100001000" => q_unbuf <= my_rom(7944);
      when "1111100001001" => q_unbuf <= my_rom(7945);
      when "1111100001010" => q_unbuf <= my_rom(7946);
      when "1111100001011" => q_unbuf <= my_rom(7947);
      when "1111100001100" => q_unbuf <= my_rom(7948);
      when "1111100001101" => q_unbuf <= my_rom(7949);
      when "1111100001110" => q_unbuf <= my_rom(7950);
      when "1111100001111" => q_unbuf <= my_rom(7951);
      when "1111100010000" => q_unbuf <= my_rom(7952);
      when "1111100010001" => q_unbuf <= my_rom(7953);
      when "1111100010010" => q_unbuf <= my_rom(7954);
      when "1111100010011" => q_unbuf <= my_rom(7955);
      when "1111100010100" => q_unbuf <= my_rom(7956);
      when "1111100010101" => q_unbuf <= my_rom(7957);
      when "1111100010110" => q_unbuf <= my_rom(7958);
      when "1111100010111" => q_unbuf <= my_rom(7959);
      when "1111100011000" => q_unbuf <= my_rom(7960);
      when "1111100011001" => q_unbuf <= my_rom(7961);
      when "1111100011010" => q_unbuf <= my_rom(7962);
      when "1111100011011" => q_unbuf <= my_rom(7963);
      when "1111100011100" => q_unbuf <= my_rom(7964);
      when "1111100011101" => q_unbuf <= my_rom(7965);
      when "1111100011110" => q_unbuf <= my_rom(7966);
      when "1111100011111" => q_unbuf <= my_rom(7967);
      when "1111100100000" => q_unbuf <= my_rom(7968);
      when "1111100100001" => q_unbuf <= my_rom(7969);
      when "1111100100010" => q_unbuf <= my_rom(7970);
      when "1111100100011" => q_unbuf <= my_rom(7971);
      when "1111100100100" => q_unbuf <= my_rom(7972);
      when "1111100100101" => q_unbuf <= my_rom(7973);
      when "1111100100110" => q_unbuf <= my_rom(7974);
      when "1111100100111" => q_unbuf <= my_rom(7975);
      when "1111100101000" => q_unbuf <= my_rom(7976);
      when "1111100101001" => q_unbuf <= my_rom(7977);
      when "1111100101010" => q_unbuf <= my_rom(7978);
      when "1111100101011" => q_unbuf <= my_rom(7979);
      when "1111100101100" => q_unbuf <= my_rom(7980);
      when "1111100101101" => q_unbuf <= my_rom(7981);
      when "1111100101110" => q_unbuf <= my_rom(7982);
      when "1111100101111" => q_unbuf <= my_rom(7983);
      when "1111100110000" => q_unbuf <= my_rom(7984);
      when "1111100110001" => q_unbuf <= my_rom(7985);
      when "1111100110010" => q_unbuf <= my_rom(7986);
      when "1111100110011" => q_unbuf <= my_rom(7987);
      when "1111100110100" => q_unbuf <= my_rom(7988);
      when "1111100110101" => q_unbuf <= my_rom(7989);
      when "1111100110110" => q_unbuf <= my_rom(7990);
      when "1111100110111" => q_unbuf <= my_rom(7991);
      when "1111100111000" => q_unbuf <= my_rom(7992);
      when "1111100111001" => q_unbuf <= my_rom(7993);
      when "1111100111010" => q_unbuf <= my_rom(7994);
      when "1111100111011" => q_unbuf <= my_rom(7995);
      when "1111100111100" => q_unbuf <= my_rom(7996);
      when "1111100111101" => q_unbuf <= my_rom(7997);
      when "1111100111110" => q_unbuf <= my_rom(7998);
      when "1111100111111" => q_unbuf <= my_rom(7999);
      when "1111101000000" => q_unbuf <= my_rom(8000);
      when "1111101000001" => q_unbuf <= my_rom(8001);
      when "1111101000010" => q_unbuf <= my_rom(8002);
      when "1111101000011" => q_unbuf <= my_rom(8003);
      when "1111101000100" => q_unbuf <= my_rom(8004);
      when "1111101000101" => q_unbuf <= my_rom(8005);
      when "1111101000110" => q_unbuf <= my_rom(8006);
      when "1111101000111" => q_unbuf <= my_rom(8007);
      when "1111101001000" => q_unbuf <= my_rom(8008);
      when "1111101001001" => q_unbuf <= my_rom(8009);
      when "1111101001010" => q_unbuf <= my_rom(8010);
      when "1111101001011" => q_unbuf <= my_rom(8011);
      when "1111101001100" => q_unbuf <= my_rom(8012);
      when "1111101001101" => q_unbuf <= my_rom(8013);
      when "1111101001110" => q_unbuf <= my_rom(8014);
      when "1111101001111" => q_unbuf <= my_rom(8015);
      when "1111101010000" => q_unbuf <= my_rom(8016);
      when "1111101010001" => q_unbuf <= my_rom(8017);
      when "1111101010010" => q_unbuf <= my_rom(8018);
      when "1111101010011" => q_unbuf <= my_rom(8019);
      when "1111101010100" => q_unbuf <= my_rom(8020);
      when "1111101010101" => q_unbuf <= my_rom(8021);
      when "1111101010110" => q_unbuf <= my_rom(8022);
      when "1111101010111" => q_unbuf <= my_rom(8023);
      when "1111101011000" => q_unbuf <= my_rom(8024);
      when "1111101011001" => q_unbuf <= my_rom(8025);
      when "1111101011010" => q_unbuf <= my_rom(8026);
      when "1111101011011" => q_unbuf <= my_rom(8027);
      when "1111101011100" => q_unbuf <= my_rom(8028);
      when "1111101011101" => q_unbuf <= my_rom(8029);
      when "1111101011110" => q_unbuf <= my_rom(8030);
      when "1111101011111" => q_unbuf <= my_rom(8031);
      when "1111101100000" => q_unbuf <= my_rom(8032);
      when "1111101100001" => q_unbuf <= my_rom(8033);
      when "1111101100010" => q_unbuf <= my_rom(8034);
      when "1111101100011" => q_unbuf <= my_rom(8035);
      when "1111101100100" => q_unbuf <= my_rom(8036);
      when "1111101100101" => q_unbuf <= my_rom(8037);
      when "1111101100110" => q_unbuf <= my_rom(8038);
      when "1111101100111" => q_unbuf <= my_rom(8039);
      when "1111101101000" => q_unbuf <= my_rom(8040);
      when "1111101101001" => q_unbuf <= my_rom(8041);
      when "1111101101010" => q_unbuf <= my_rom(8042);
      when "1111101101011" => q_unbuf <= my_rom(8043);
      when "1111101101100" => q_unbuf <= my_rom(8044);
      when "1111101101101" => q_unbuf <= my_rom(8045);
      when "1111101101110" => q_unbuf <= my_rom(8046);
      when "1111101101111" => q_unbuf <= my_rom(8047);
      when "1111101110000" => q_unbuf <= my_rom(8048);
      when "1111101110001" => q_unbuf <= my_rom(8049);
      when "1111101110010" => q_unbuf <= my_rom(8050);
      when "1111101110011" => q_unbuf <= my_rom(8051);
      when "1111101110100" => q_unbuf <= my_rom(8052);
      when "1111101110101" => q_unbuf <= my_rom(8053);
      when "1111101110110" => q_unbuf <= my_rom(8054);
      when "1111101110111" => q_unbuf <= my_rom(8055);
      when "1111101111000" => q_unbuf <= my_rom(8056);
      when "1111101111001" => q_unbuf <= my_rom(8057);
      when "1111101111010" => q_unbuf <= my_rom(8058);
      when "1111101111011" => q_unbuf <= my_rom(8059);
      when "1111101111100" => q_unbuf <= my_rom(8060);
      when "1111101111101" => q_unbuf <= my_rom(8061);
      when "1111101111110" => q_unbuf <= my_rom(8062);
      when "1111101111111" => q_unbuf <= my_rom(8063);
      when "1111110000000" => q_unbuf <= my_rom(8064);
      when "1111110000001" => q_unbuf <= my_rom(8065);
      when "1111110000010" => q_unbuf <= my_rom(8066);
      when "1111110000011" => q_unbuf <= my_rom(8067);
      when "1111110000100" => q_unbuf <= my_rom(8068);
      when "1111110000101" => q_unbuf <= my_rom(8069);
      when "1111110000110" => q_unbuf <= my_rom(8070);
      when "1111110000111" => q_unbuf <= my_rom(8071);
      when "1111110001000" => q_unbuf <= my_rom(8072);
      when "1111110001001" => q_unbuf <= my_rom(8073);
      when "1111110001010" => q_unbuf <= my_rom(8074);
      when "1111110001011" => q_unbuf <= my_rom(8075);
      when "1111110001100" => q_unbuf <= my_rom(8076);
      when "1111110001101" => q_unbuf <= my_rom(8077);
      when "1111110001110" => q_unbuf <= my_rom(8078);
      when "1111110001111" => q_unbuf <= my_rom(8079);
      when "1111110010000" => q_unbuf <= my_rom(8080);
      when "1111110010001" => q_unbuf <= my_rom(8081);
      when "1111110010010" => q_unbuf <= my_rom(8082);
      when "1111110010011" => q_unbuf <= my_rom(8083);
      when "1111110010100" => q_unbuf <= my_rom(8084);
      when "1111110010101" => q_unbuf <= my_rom(8085);
      when "1111110010110" => q_unbuf <= my_rom(8086);
      when "1111110010111" => q_unbuf <= my_rom(8087);
      when "1111110011000" => q_unbuf <= my_rom(8088);
      when "1111110011001" => q_unbuf <= my_rom(8089);
      when "1111110011010" => q_unbuf <= my_rom(8090);
      when "1111110011011" => q_unbuf <= my_rom(8091);
      when "1111110011100" => q_unbuf <= my_rom(8092);
      when "1111110011101" => q_unbuf <= my_rom(8093);
      when "1111110011110" => q_unbuf <= my_rom(8094);
      when "1111110011111" => q_unbuf <= my_rom(8095);
      when "1111110100000" => q_unbuf <= my_rom(8096);
      when "1111110100001" => q_unbuf <= my_rom(8097);
      when "1111110100010" => q_unbuf <= my_rom(8098);
      when "1111110100011" => q_unbuf <= my_rom(8099);
      when "1111110100100" => q_unbuf <= my_rom(8100);
      when "1111110100101" => q_unbuf <= my_rom(8101);
      when "1111110100110" => q_unbuf <= my_rom(8102);
      when "1111110100111" => q_unbuf <= my_rom(8103);
      when "1111110101000" => q_unbuf <= my_rom(8104);
      when "1111110101001" => q_unbuf <= my_rom(8105);
      when "1111110101010" => q_unbuf <= my_rom(8106);
      when "1111110101011" => q_unbuf <= my_rom(8107);
      when "1111110101100" => q_unbuf <= my_rom(8108);
      when "1111110101101" => q_unbuf <= my_rom(8109);
      when "1111110101110" => q_unbuf <= my_rom(8110);
      when "1111110101111" => q_unbuf <= my_rom(8111);
      when "1111110110000" => q_unbuf <= my_rom(8112);
      when "1111110110001" => q_unbuf <= my_rom(8113);
      when "1111110110010" => q_unbuf <= my_rom(8114);
      when "1111110110011" => q_unbuf <= my_rom(8115);
      when "1111110110100" => q_unbuf <= my_rom(8116);
      when "1111110110101" => q_unbuf <= my_rom(8117);
      when "1111110110110" => q_unbuf <= my_rom(8118);
      when "1111110110111" => q_unbuf <= my_rom(8119);
      when "1111110111000" => q_unbuf <= my_rom(8120);
      when "1111110111001" => q_unbuf <= my_rom(8121);
      when "1111110111010" => q_unbuf <= my_rom(8122);
      when "1111110111011" => q_unbuf <= my_rom(8123);
      when "1111110111100" => q_unbuf <= my_rom(8124);
      when "1111110111101" => q_unbuf <= my_rom(8125);
      when "1111110111110" => q_unbuf <= my_rom(8126);
      when "1111110111111" => q_unbuf <= my_rom(8127);
      when "1111111000000" => q_unbuf <= my_rom(8128);
      when "1111111000001" => q_unbuf <= my_rom(8129);
      when "1111111000010" => q_unbuf <= my_rom(8130);
      when "1111111000011" => q_unbuf <= my_rom(8131);
      when "1111111000100" => q_unbuf <= my_rom(8132);
      when "1111111000101" => q_unbuf <= my_rom(8133);
      when "1111111000110" => q_unbuf <= my_rom(8134);
      when "1111111000111" => q_unbuf <= my_rom(8135);
      when "1111111001000" => q_unbuf <= my_rom(8136);
      when "1111111001001" => q_unbuf <= my_rom(8137);
      when "1111111001010" => q_unbuf <= my_rom(8138);
      when "1111111001011" => q_unbuf <= my_rom(8139);
      when "1111111001100" => q_unbuf <= my_rom(8140);
      when "1111111001101" => q_unbuf <= my_rom(8141);
      when "1111111001110" => q_unbuf <= my_rom(8142);
      when "1111111001111" => q_unbuf <= my_rom(8143);
      when "1111111010000" => q_unbuf <= my_rom(8144);
      when "1111111010001" => q_unbuf <= my_rom(8145);
      when "1111111010010" => q_unbuf <= my_rom(8146);
      when "1111111010011" => q_unbuf <= my_rom(8147);
      when "1111111010100" => q_unbuf <= my_rom(8148);
      when "1111111010101" => q_unbuf <= my_rom(8149);
      when "1111111010110" => q_unbuf <= my_rom(8150);
      when "1111111010111" => q_unbuf <= my_rom(8151);
      when "1111111011000" => q_unbuf <= my_rom(8152);
      when "1111111011001" => q_unbuf <= my_rom(8153);
      when "1111111011010" => q_unbuf <= my_rom(8154);
      when "1111111011011" => q_unbuf <= my_rom(8155);
      when "1111111011100" => q_unbuf <= my_rom(8156);
      when "1111111011101" => q_unbuf <= my_rom(8157);
      when "1111111011110" => q_unbuf <= my_rom(8158);
      when "1111111011111" => q_unbuf <= my_rom(8159);
      when "1111111100000" => q_unbuf <= my_rom(8160);
      when "1111111100001" => q_unbuf <= my_rom(8161);
      when "1111111100010" => q_unbuf <= my_rom(8162);
      when "1111111100011" => q_unbuf <= my_rom(8163);
      when "1111111100100" => q_unbuf <= my_rom(8164);
      when "1111111100101" => q_unbuf <= my_rom(8165);
      when "1111111100110" => q_unbuf <= my_rom(8166);
      when "1111111100111" => q_unbuf <= my_rom(8167);
      when "1111111101000" => q_unbuf <= my_rom(8168);
      when "1111111101001" => q_unbuf <= my_rom(8169);
      when "1111111101010" => q_unbuf <= my_rom(8170);
      when "1111111101011" => q_unbuf <= my_rom(8171);
      when "1111111101100" => q_unbuf <= my_rom(8172);
      when "1111111101101" => q_unbuf <= my_rom(8173);
      when "1111111101110" => q_unbuf <= my_rom(8174);
      when "1111111101111" => q_unbuf <= my_rom(8175);
      when "1111111110000" => q_unbuf <= my_rom(8176);
      when "1111111110001" => q_unbuf <= my_rom(8177);
      when "1111111110010" => q_unbuf <= my_rom(8178);
      when "1111111110011" => q_unbuf <= my_rom(8179);
      when "1111111110100" => q_unbuf <= my_rom(8180);
      when "1111111110101" => q_unbuf <= my_rom(8181);
      when "1111111110110" => q_unbuf <= my_rom(8182);
      when "1111111110111" => q_unbuf <= my_rom(8183);
      when "1111111111000" => q_unbuf <= my_rom(8184);
      when "1111111111001" => q_unbuf <= my_rom(8185);
      when "1111111111010" => q_unbuf <= my_rom(8186);
      when "1111111111011" => q_unbuf <= my_rom(8187);
      when "1111111111100" => q_unbuf <= my_rom(8188);
      when "1111111111101" => q_unbuf <= my_rom(8189);
      when "1111111111110" => q_unbuf <= my_rom(8190);
      when "1111111111111" => q_unbuf <= my_rom(8191);
      when others => q_unbuf <= "00000000";
     end case;
  end process;

  process
  begin
    wait until rising_edge(clock);
    q <= q_unbuf;
  end process;

end architecture behavioral;
